
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"00",x"00",x"18",x"3c"),
     1 => (x"24",x"24",x"3c",x"18"),
     2 => (x"00",x"00",x"fc",x"fc"),
     3 => (x"04",x"04",x"7c",x"7c"),
     4 => (x"00",x"00",x"08",x"0c"),
     5 => (x"54",x"54",x"5c",x"48"),
     6 => (x"00",x"00",x"20",x"74"),
     7 => (x"44",x"7f",x"3f",x"04"),
     8 => (x"00",x"00",x"00",x"44"),
     9 => (x"40",x"40",x"7c",x"3c"),
    10 => (x"00",x"00",x"7c",x"7c"),
    11 => (x"60",x"60",x"3c",x"1c"),
    12 => (x"3c",x"00",x"1c",x"3c"),
    13 => (x"60",x"30",x"60",x"7c"),
    14 => (x"44",x"00",x"3c",x"7c"),
    15 => (x"38",x"10",x"38",x"6c"),
    16 => (x"00",x"00",x"44",x"6c"),
    17 => (x"60",x"e0",x"bc",x"1c"),
    18 => (x"00",x"00",x"1c",x"3c"),
    19 => (x"5c",x"74",x"64",x"44"),
    20 => (x"00",x"00",x"44",x"4c"),
    21 => (x"77",x"3e",x"08",x"08"),
    22 => (x"00",x"00",x"41",x"41"),
    23 => (x"7f",x"7f",x"00",x"00"),
    24 => (x"00",x"00",x"00",x"00"),
    25 => (x"3e",x"77",x"41",x"41"),
    26 => (x"02",x"00",x"08",x"08"),
    27 => (x"02",x"03",x"01",x"01"),
    28 => (x"7f",x"00",x"01",x"02"),
    29 => (x"7f",x"7f",x"7f",x"7f"),
    30 => (x"08",x"00",x"7f",x"7f"),
    31 => (x"3e",x"1c",x"1c",x"08"),
    32 => (x"7f",x"7f",x"7f",x"3e"),
    33 => (x"1c",x"3e",x"3e",x"7f"),
    34 => (x"00",x"08",x"08",x"1c"),
    35 => (x"7c",x"7c",x"18",x"10"),
    36 => (x"00",x"00",x"10",x"18"),
    37 => (x"7c",x"7c",x"30",x"10"),
    38 => (x"10",x"00",x"10",x"30"),
    39 => (x"78",x"60",x"60",x"30"),
    40 => (x"42",x"00",x"06",x"1e"),
    41 => (x"3c",x"18",x"3c",x"66"),
    42 => (x"78",x"00",x"42",x"66"),
    43 => (x"c6",x"c2",x"6a",x"38"),
    44 => (x"60",x"00",x"38",x"6c"),
    45 => (x"00",x"60",x"00",x"00"),
    46 => (x"0e",x"00",x"60",x"00"),
    47 => (x"5d",x"5c",x"5b",x"5e"),
    48 => (x"4c",x"71",x"1e",x"0e"),
    49 => (x"bf",x"d9",x"ec",x"c2"),
    50 => (x"c0",x"4b",x"c0",x"4d"),
    51 => (x"02",x"ab",x"74",x"1e"),
    52 => (x"a6",x"c4",x"87",x"c7"),
    53 => (x"c5",x"78",x"c0",x"48"),
    54 => (x"48",x"a6",x"c4",x"87"),
    55 => (x"66",x"c4",x"78",x"c1"),
    56 => (x"ee",x"49",x"73",x"1e"),
    57 => (x"86",x"c8",x"87",x"df"),
    58 => (x"ef",x"49",x"e0",x"c0"),
    59 => (x"a5",x"c4",x"87",x"ee"),
    60 => (x"f0",x"49",x"6a",x"4a"),
    61 => (x"c6",x"f1",x"87",x"f0"),
    62 => (x"c1",x"85",x"cb",x"87"),
    63 => (x"ab",x"b7",x"c8",x"83"),
    64 => (x"87",x"c7",x"ff",x"04"),
    65 => (x"26",x"4d",x"26",x"26"),
    66 => (x"26",x"4b",x"26",x"4c"),
    67 => (x"4a",x"71",x"1e",x"4f"),
    68 => (x"5a",x"dd",x"ec",x"c2"),
    69 => (x"48",x"dd",x"ec",x"c2"),
    70 => (x"fe",x"49",x"78",x"c7"),
    71 => (x"4f",x"26",x"87",x"dd"),
    72 => (x"71",x"1e",x"73",x"1e"),
    73 => (x"aa",x"b7",x"c0",x"4a"),
    74 => (x"c2",x"87",x"d3",x"03"),
    75 => (x"05",x"bf",x"dc",x"d2"),
    76 => (x"4b",x"c1",x"87",x"c4"),
    77 => (x"4b",x"c0",x"87",x"c2"),
    78 => (x"5b",x"e0",x"d2",x"c2"),
    79 => (x"d2",x"c2",x"87",x"c4"),
    80 => (x"d2",x"c2",x"5a",x"e0"),
    81 => (x"c1",x"4a",x"bf",x"dc"),
    82 => (x"a2",x"c0",x"c1",x"9a"),
    83 => (x"87",x"e8",x"ec",x"49"),
    84 => (x"d2",x"c2",x"48",x"fc"),
    85 => (x"fe",x"78",x"bf",x"dc"),
    86 => (x"71",x"1e",x"87",x"ef"),
    87 => (x"1e",x"66",x"c4",x"4a"),
    88 => (x"f9",x"ea",x"49",x"72"),
    89 => (x"4f",x"26",x"26",x"87"),
    90 => (x"48",x"d4",x"ff",x"1e"),
    91 => (x"ff",x"78",x"ff",x"c3"),
    92 => (x"e1",x"c0",x"48",x"d0"),
    93 => (x"48",x"d4",x"ff",x"78"),
    94 => (x"48",x"71",x"78",x"c1"),
    95 => (x"d4",x"ff",x"30",x"c4"),
    96 => (x"d0",x"ff",x"78",x"08"),
    97 => (x"78",x"e0",x"c0",x"48"),
    98 => (x"c2",x"1e",x"4f",x"26"),
    99 => (x"49",x"bf",x"dc",x"d2"),
   100 => (x"c2",x"87",x"f9",x"e6"),
   101 => (x"e8",x"48",x"d1",x"ec"),
   102 => (x"ec",x"c2",x"78",x"bf"),
   103 => (x"bf",x"ec",x"48",x"cd"),
   104 => (x"d1",x"ec",x"c2",x"78"),
   105 => (x"c3",x"49",x"4a",x"bf"),
   106 => (x"b7",x"c8",x"99",x"ff"),
   107 => (x"71",x"48",x"72",x"2a"),
   108 => (x"d9",x"ec",x"c2",x"b0"),
   109 => (x"0e",x"4f",x"26",x"58"),
   110 => (x"5d",x"5c",x"5b",x"5e"),
   111 => (x"ff",x"4b",x"71",x"0e"),
   112 => (x"ec",x"c2",x"87",x"c8"),
   113 => (x"50",x"c0",x"48",x"cc"),
   114 => (x"df",x"e6",x"49",x"73"),
   115 => (x"4c",x"49",x"70",x"87"),
   116 => (x"ee",x"cb",x"9c",x"c2"),
   117 => (x"87",x"cc",x"cb",x"49"),
   118 => (x"ec",x"c2",x"4d",x"70"),
   119 => (x"05",x"bf",x"97",x"cc"),
   120 => (x"d0",x"87",x"e2",x"c1"),
   121 => (x"ec",x"c2",x"49",x"66"),
   122 => (x"05",x"99",x"bf",x"d5"),
   123 => (x"66",x"d4",x"87",x"d6"),
   124 => (x"cd",x"ec",x"c2",x"49"),
   125 => (x"cb",x"05",x"99",x"bf"),
   126 => (x"e5",x"49",x"73",x"87"),
   127 => (x"98",x"70",x"87",x"ee"),
   128 => (x"87",x"c1",x"c1",x"02"),
   129 => (x"c1",x"fe",x"4c",x"c1"),
   130 => (x"ca",x"49",x"75",x"87"),
   131 => (x"98",x"70",x"87",x"e2"),
   132 => (x"c2",x"87",x"c6",x"02"),
   133 => (x"c1",x"48",x"cc",x"ec"),
   134 => (x"cc",x"ec",x"c2",x"50"),
   135 => (x"c0",x"05",x"bf",x"97"),
   136 => (x"ec",x"c2",x"87",x"e3"),
   137 => (x"d0",x"49",x"bf",x"d5"),
   138 => (x"ff",x"05",x"99",x"66"),
   139 => (x"ec",x"c2",x"87",x"d6"),
   140 => (x"d4",x"49",x"bf",x"cd"),
   141 => (x"ff",x"05",x"99",x"66"),
   142 => (x"49",x"73",x"87",x"ca"),
   143 => (x"70",x"87",x"ed",x"e4"),
   144 => (x"ff",x"fe",x"05",x"98"),
   145 => (x"fa",x"48",x"74",x"87"),
   146 => (x"5e",x"0e",x"87",x"fb"),
   147 => (x"0e",x"5d",x"5c",x"5b"),
   148 => (x"4d",x"c0",x"86",x"f8"),
   149 => (x"7e",x"bf",x"ec",x"4c"),
   150 => (x"c2",x"48",x"a6",x"c4"),
   151 => (x"78",x"bf",x"d9",x"ec"),
   152 => (x"1e",x"c0",x"1e",x"c1"),
   153 => (x"ce",x"fd",x"49",x"c7"),
   154 => (x"70",x"86",x"c8",x"87"),
   155 => (x"87",x"cd",x"02",x"98"),
   156 => (x"eb",x"fa",x"49",x"ff"),
   157 => (x"49",x"da",x"c1",x"87"),
   158 => (x"c1",x"87",x"f1",x"e3"),
   159 => (x"cc",x"ec",x"c2",x"4d"),
   160 => (x"cf",x"02",x"bf",x"97"),
   161 => (x"d4",x"d2",x"c2",x"87"),
   162 => (x"b9",x"c1",x"49",x"bf"),
   163 => (x"59",x"d8",x"d2",x"c2"),
   164 => (x"87",x"d4",x"fb",x"71"),
   165 => (x"bf",x"d1",x"ec",x"c2"),
   166 => (x"dc",x"d2",x"c2",x"4b"),
   167 => (x"e9",x"c0",x"05",x"bf"),
   168 => (x"49",x"fd",x"c3",x"87"),
   169 => (x"c3",x"87",x"c5",x"e3"),
   170 => (x"ff",x"e2",x"49",x"fa"),
   171 => (x"c3",x"49",x"73",x"87"),
   172 => (x"1e",x"71",x"99",x"ff"),
   173 => (x"e1",x"fa",x"49",x"c0"),
   174 => (x"c8",x"49",x"73",x"87"),
   175 => (x"1e",x"71",x"29",x"b7"),
   176 => (x"d5",x"fa",x"49",x"c1"),
   177 => (x"c5",x"86",x"c8",x"87"),
   178 => (x"ec",x"c2",x"87",x"f4"),
   179 => (x"9b",x"4b",x"bf",x"d5"),
   180 => (x"c2",x"87",x"dd",x"02"),
   181 => (x"49",x"bf",x"d8",x"d2"),
   182 => (x"70",x"87",x"d5",x"c7"),
   183 => (x"87",x"c4",x"05",x"98"),
   184 => (x"87",x"d2",x"4b",x"c0"),
   185 => (x"c6",x"49",x"e0",x"c2"),
   186 => (x"d2",x"c2",x"87",x"fa"),
   187 => (x"87",x"c6",x"58",x"dc"),
   188 => (x"48",x"d8",x"d2",x"c2"),
   189 => (x"49",x"73",x"78",x"c0"),
   190 => (x"cd",x"05",x"99",x"c2"),
   191 => (x"49",x"eb",x"c3",x"87"),
   192 => (x"70",x"87",x"e9",x"e1"),
   193 => (x"02",x"99",x"c2",x"49"),
   194 => (x"4c",x"fb",x"87",x"c2"),
   195 => (x"99",x"c1",x"49",x"73"),
   196 => (x"c3",x"87",x"cd",x"05"),
   197 => (x"d3",x"e1",x"49",x"f4"),
   198 => (x"c2",x"49",x"70",x"87"),
   199 => (x"87",x"c2",x"02",x"99"),
   200 => (x"49",x"73",x"4c",x"fa"),
   201 => (x"cd",x"05",x"99",x"c8"),
   202 => (x"49",x"f5",x"c3",x"87"),
   203 => (x"70",x"87",x"fd",x"e0"),
   204 => (x"02",x"99",x"c2",x"49"),
   205 => (x"ec",x"c2",x"87",x"d5"),
   206 => (x"ca",x"02",x"bf",x"dd"),
   207 => (x"88",x"c1",x"48",x"87"),
   208 => (x"58",x"e1",x"ec",x"c2"),
   209 => (x"ff",x"87",x"c2",x"c0"),
   210 => (x"73",x"4d",x"c1",x"4c"),
   211 => (x"05",x"99",x"c4",x"49"),
   212 => (x"f2",x"c3",x"87",x"cd"),
   213 => (x"87",x"d4",x"e0",x"49"),
   214 => (x"99",x"c2",x"49",x"70"),
   215 => (x"c2",x"87",x"dc",x"02"),
   216 => (x"7e",x"bf",x"dd",x"ec"),
   217 => (x"a8",x"b7",x"c7",x"48"),
   218 => (x"87",x"cb",x"c0",x"03"),
   219 => (x"80",x"c1",x"48",x"6e"),
   220 => (x"58",x"e1",x"ec",x"c2"),
   221 => (x"fe",x"87",x"c2",x"c0"),
   222 => (x"c3",x"4d",x"c1",x"4c"),
   223 => (x"df",x"ff",x"49",x"fd"),
   224 => (x"49",x"70",x"87",x"ea"),
   225 => (x"d5",x"02",x"99",x"c2"),
   226 => (x"dd",x"ec",x"c2",x"87"),
   227 => (x"c9",x"c0",x"02",x"bf"),
   228 => (x"dd",x"ec",x"c2",x"87"),
   229 => (x"c0",x"78",x"c0",x"48"),
   230 => (x"4c",x"fd",x"87",x"c2"),
   231 => (x"fa",x"c3",x"4d",x"c1"),
   232 => (x"c7",x"df",x"ff",x"49"),
   233 => (x"c2",x"49",x"70",x"87"),
   234 => (x"d9",x"c0",x"02",x"99"),
   235 => (x"dd",x"ec",x"c2",x"87"),
   236 => (x"b7",x"c7",x"48",x"bf"),
   237 => (x"c9",x"c0",x"03",x"a8"),
   238 => (x"dd",x"ec",x"c2",x"87"),
   239 => (x"c0",x"78",x"c7",x"48"),
   240 => (x"4c",x"fc",x"87",x"c2"),
   241 => (x"b7",x"c0",x"4d",x"c1"),
   242 => (x"d3",x"c0",x"03",x"ac"),
   243 => (x"48",x"66",x"c4",x"87"),
   244 => (x"70",x"80",x"d8",x"c1"),
   245 => (x"02",x"bf",x"6e",x"7e"),
   246 => (x"4b",x"87",x"c5",x"c0"),
   247 => (x"0f",x"73",x"49",x"74"),
   248 => (x"f0",x"c3",x"1e",x"c0"),
   249 => (x"49",x"da",x"c1",x"1e"),
   250 => (x"c8",x"87",x"cc",x"f7"),
   251 => (x"02",x"98",x"70",x"86"),
   252 => (x"c2",x"87",x"d8",x"c0"),
   253 => (x"7e",x"bf",x"dd",x"ec"),
   254 => (x"91",x"cb",x"49",x"6e"),
   255 => (x"71",x"4a",x"66",x"c4"),
   256 => (x"c0",x"02",x"6a",x"82"),
   257 => (x"6e",x"4b",x"87",x"c5"),
   258 => (x"75",x"0f",x"73",x"49"),
   259 => (x"c8",x"c0",x"02",x"9d"),
   260 => (x"dd",x"ec",x"c2",x"87"),
   261 => (x"e2",x"f2",x"49",x"bf"),
   262 => (x"e0",x"d2",x"c2",x"87"),
   263 => (x"dd",x"c0",x"02",x"bf"),
   264 => (x"cb",x"c2",x"49",x"87"),
   265 => (x"02",x"98",x"70",x"87"),
   266 => (x"c2",x"87",x"d3",x"c0"),
   267 => (x"49",x"bf",x"dd",x"ec"),
   268 => (x"c0",x"87",x"c8",x"f2"),
   269 => (x"87",x"e8",x"f3",x"49"),
   270 => (x"48",x"e0",x"d2",x"c2"),
   271 => (x"8e",x"f8",x"78",x"c0"),
   272 => (x"0e",x"87",x"c2",x"f3"),
   273 => (x"5d",x"5c",x"5b",x"5e"),
   274 => (x"4c",x"71",x"1e",x"0e"),
   275 => (x"bf",x"d9",x"ec",x"c2"),
   276 => (x"a1",x"cd",x"c1",x"49"),
   277 => (x"81",x"d1",x"c1",x"4d"),
   278 => (x"9c",x"74",x"7e",x"69"),
   279 => (x"c4",x"87",x"cf",x"02"),
   280 => (x"7b",x"74",x"4b",x"a5"),
   281 => (x"bf",x"d9",x"ec",x"c2"),
   282 => (x"87",x"e1",x"f2",x"49"),
   283 => (x"9c",x"74",x"7b",x"6e"),
   284 => (x"c0",x"87",x"c4",x"05"),
   285 => (x"c1",x"87",x"c2",x"4b"),
   286 => (x"f2",x"49",x"73",x"4b"),
   287 => (x"66",x"d4",x"87",x"e2"),
   288 => (x"49",x"87",x"c7",x"02"),
   289 => (x"4a",x"70",x"87",x"de"),
   290 => (x"4a",x"c0",x"87",x"c2"),
   291 => (x"5a",x"e4",x"d2",x"c2"),
   292 => (x"87",x"f1",x"f1",x"26"),
   293 => (x"00",x"00",x"00",x"00"),
   294 => (x"00",x"00",x"00",x"00"),
   295 => (x"00",x"00",x"00",x"00"),
   296 => (x"00",x"00",x"00",x"00"),
   297 => (x"ff",x"4a",x"71",x"1e"),
   298 => (x"72",x"49",x"bf",x"c8"),
   299 => (x"4f",x"26",x"48",x"a1"),
   300 => (x"bf",x"c8",x"ff",x"1e"),
   301 => (x"c0",x"c0",x"fe",x"89"),
   302 => (x"a9",x"c0",x"c0",x"c0"),
   303 => (x"c0",x"87",x"c4",x"01"),
   304 => (x"c1",x"87",x"c2",x"4a"),
   305 => (x"26",x"48",x"72",x"4a"),
   306 => (x"5b",x"5e",x"0e",x"4f"),
   307 => (x"71",x"0e",x"5d",x"5c"),
   308 => (x"4c",x"d4",x"ff",x"4b"),
   309 => (x"c0",x"48",x"66",x"d0"),
   310 => (x"ff",x"49",x"d6",x"78"),
   311 => (x"c3",x"87",x"c5",x"dc"),
   312 => (x"49",x"6c",x"7c",x"ff"),
   313 => (x"71",x"99",x"ff",x"c3"),
   314 => (x"f0",x"c3",x"49",x"4d"),
   315 => (x"a9",x"e0",x"c1",x"99"),
   316 => (x"c3",x"87",x"cb",x"05"),
   317 => (x"48",x"6c",x"7c",x"ff"),
   318 => (x"66",x"d0",x"98",x"c3"),
   319 => (x"ff",x"c3",x"78",x"08"),
   320 => (x"49",x"4a",x"6c",x"7c"),
   321 => (x"ff",x"c3",x"31",x"c8"),
   322 => (x"71",x"4a",x"6c",x"7c"),
   323 => (x"c8",x"49",x"72",x"b2"),
   324 => (x"7c",x"ff",x"c3",x"31"),
   325 => (x"b2",x"71",x"4a",x"6c"),
   326 => (x"31",x"c8",x"49",x"72"),
   327 => (x"6c",x"7c",x"ff",x"c3"),
   328 => (x"ff",x"b2",x"71",x"4a"),
   329 => (x"e0",x"c0",x"48",x"d0"),
   330 => (x"02",x"9b",x"73",x"78"),
   331 => (x"7b",x"72",x"87",x"c2"),
   332 => (x"4d",x"26",x"48",x"75"),
   333 => (x"4b",x"26",x"4c",x"26"),
   334 => (x"26",x"1e",x"4f",x"26"),
   335 => (x"5b",x"5e",x"0e",x"4f"),
   336 => (x"86",x"f8",x"0e",x"5c"),
   337 => (x"a6",x"c8",x"1e",x"76"),
   338 => (x"87",x"fd",x"fd",x"49"),
   339 => (x"4b",x"70",x"86",x"c4"),
   340 => (x"a8",x"c8",x"48",x"6e"),
   341 => (x"87",x"f0",x"c2",x"03"),
   342 => (x"f0",x"c3",x"4a",x"73"),
   343 => (x"aa",x"d0",x"c1",x"9a"),
   344 => (x"c1",x"87",x"c7",x"02"),
   345 => (x"c2",x"05",x"aa",x"e0"),
   346 => (x"49",x"73",x"87",x"de"),
   347 => (x"c3",x"02",x"99",x"c8"),
   348 => (x"87",x"c6",x"ff",x"87"),
   349 => (x"9c",x"c3",x"4c",x"73"),
   350 => (x"c1",x"05",x"ac",x"c2"),
   351 => (x"66",x"c4",x"87",x"c2"),
   352 => (x"71",x"31",x"c9",x"49"),
   353 => (x"4a",x"66",x"c4",x"1e"),
   354 => (x"ec",x"c2",x"92",x"d4"),
   355 => (x"81",x"72",x"49",x"e1"),
   356 => (x"87",x"f3",x"d0",x"fe"),
   357 => (x"d9",x"ff",x"49",x"d8"),
   358 => (x"c0",x"c8",x"87",x"ca"),
   359 => (x"fe",x"da",x"c2",x"1e"),
   360 => (x"f9",x"ec",x"fd",x"49"),
   361 => (x"48",x"d0",x"ff",x"87"),
   362 => (x"c2",x"78",x"e0",x"c0"),
   363 => (x"cc",x"1e",x"fe",x"da"),
   364 => (x"92",x"d4",x"4a",x"66"),
   365 => (x"49",x"e1",x"ec",x"c2"),
   366 => (x"ce",x"fe",x"81",x"72"),
   367 => (x"86",x"cc",x"87",x"fb"),
   368 => (x"c1",x"05",x"ac",x"c1"),
   369 => (x"66",x"c4",x"87",x"c2"),
   370 => (x"71",x"31",x"c9",x"49"),
   371 => (x"4a",x"66",x"c4",x"1e"),
   372 => (x"ec",x"c2",x"92",x"d4"),
   373 => (x"81",x"72",x"49",x"e1"),
   374 => (x"87",x"eb",x"cf",x"fe"),
   375 => (x"1e",x"fe",x"da",x"c2"),
   376 => (x"d4",x"4a",x"66",x"c8"),
   377 => (x"e1",x"ec",x"c2",x"92"),
   378 => (x"fe",x"81",x"72",x"49"),
   379 => (x"d7",x"87",x"fc",x"cc"),
   380 => (x"ef",x"d7",x"ff",x"49"),
   381 => (x"1e",x"c0",x"c8",x"87"),
   382 => (x"49",x"fe",x"da",x"c2"),
   383 => (x"87",x"f7",x"ea",x"fd"),
   384 => (x"d0",x"ff",x"86",x"cc"),
   385 => (x"78",x"e0",x"c0",x"48"),
   386 => (x"e7",x"fc",x"8e",x"f8"),
   387 => (x"5b",x"5e",x"0e",x"87"),
   388 => (x"1e",x"0e",x"5d",x"5c"),
   389 => (x"d4",x"ff",x"4d",x"71"),
   390 => (x"7e",x"66",x"d4",x"4c"),
   391 => (x"a8",x"b7",x"c3",x"48"),
   392 => (x"c0",x"87",x"c5",x"06"),
   393 => (x"87",x"e9",x"c1",x"48"),
   394 => (x"dd",x"fe",x"49",x"75"),
   395 => (x"1e",x"75",x"87",x"e0"),
   396 => (x"d4",x"4b",x"66",x"c4"),
   397 => (x"e1",x"ec",x"c2",x"93"),
   398 => (x"fe",x"49",x"73",x"83"),
   399 => (x"c8",x"87",x"fa",x"c6"),
   400 => (x"ff",x"4b",x"6b",x"83"),
   401 => (x"e1",x"c8",x"48",x"d0"),
   402 => (x"73",x"7c",x"dd",x"78"),
   403 => (x"98",x"ff",x"c3",x"48"),
   404 => (x"49",x"73",x"7c",x"70"),
   405 => (x"71",x"29",x"b7",x"c8"),
   406 => (x"98",x"ff",x"c3",x"48"),
   407 => (x"49",x"73",x"7c",x"70"),
   408 => (x"71",x"29",x"b7",x"d0"),
   409 => (x"98",x"ff",x"c3",x"48"),
   410 => (x"48",x"73",x"7c",x"70"),
   411 => (x"70",x"28",x"b7",x"d8"),
   412 => (x"7c",x"7c",x"c0",x"7c"),
   413 => (x"7c",x"7c",x"7c",x"7c"),
   414 => (x"7c",x"7c",x"7c",x"7c"),
   415 => (x"d0",x"ff",x"7c",x"7c"),
   416 => (x"78",x"e0",x"c0",x"48"),
   417 => (x"dc",x"1e",x"66",x"c4"),
   418 => (x"fc",x"d5",x"ff",x"49"),
   419 => (x"73",x"86",x"c8",x"87"),
   420 => (x"dd",x"fa",x"26",x"48"),
   421 => (x"dd",x"fa",x"26",x"87"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

