library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c4efc287",
    12 => x"86c0c84e",
    13 => x"49c4efc2",
    14 => x"48d8dac2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087cde2",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"66c44a71",
    47 => x"88c14849",
    48 => x"7158a6c8",
    49 => x"87d40299",
    50 => x"d4ff4812",
    51 => x"66c47808",
    52 => x"88c14849",
    53 => x"7158a6c8",
    54 => x"87ec0599",
    55 => x"711e4f26",
    56 => x"4966c44a",
    57 => x"c888c148",
    58 => x"997158a6",
    59 => x"ff87d602",
    60 => x"ffc348d4",
    61 => x"c4526878",
    62 => x"c1484966",
    63 => x"58a6c888",
    64 => x"ea059971",
    65 => x"1e4f2687",
    66 => x"d4ff1e73",
    67 => x"7bffc34b",
    68 => x"ffc34a6b",
    69 => x"c8496b7b",
    70 => x"c3b17232",
    71 => x"4a6b7bff",
    72 => x"b27131c8",
    73 => x"6b7bffc3",
    74 => x"7232c849",
    75 => x"c44871b1",
    76 => x"264d2687",
    77 => x"264b264c",
    78 => x"5b5e0e4f",
    79 => x"710e5d5c",
    80 => x"4cd4ff4a",
    81 => x"ffc34872",
    82 => x"c27c7098",
    83 => x"05bfd8da",
    84 => x"66d087c8",
    85 => x"d430c948",
    86 => x"66d058a6",
    87 => x"7129d849",
    88 => x"98ffc348",
    89 => x"66d07c70",
    90 => x"7129d049",
    91 => x"98ffc348",
    92 => x"66d07c70",
    93 => x"7129c849",
    94 => x"98ffc348",
    95 => x"66d07c70",
    96 => x"98ffc348",
    97 => x"49727c70",
    98 => x"487129d0",
    99 => x"7098ffc3",
   100 => x"c94b6c7c",
   101 => x"c34dfff0",
   102 => x"d005abff",
   103 => x"7cffc387",
   104 => x"8dc14b6c",
   105 => x"c387c602",
   106 => x"f002abff",
   107 => x"fd487387",
   108 => x"c01e87ff",
   109 => x"48d4ff49",
   110 => x"c178ffc3",
   111 => x"b7c8c381",
   112 => x"87f104a9",
   113 => x"731e4f26",
   114 => x"c487e71e",
   115 => x"c04bdff8",
   116 => x"f0ffc01e",
   117 => x"fd49f7c1",
   118 => x"86c487df",
   119 => x"c005a8c1",
   120 => x"d4ff87ea",
   121 => x"78ffc348",
   122 => x"c0c0c0c1",
   123 => x"c01ec0c0",
   124 => x"e9c1f0e1",
   125 => x"87c1fd49",
   126 => x"987086c4",
   127 => x"ff87ca05",
   128 => x"ffc348d4",
   129 => x"cb48c178",
   130 => x"87e6fe87",
   131 => x"fe058bc1",
   132 => x"48c087fd",
   133 => x"1e87defc",
   134 => x"d4ff1e73",
   135 => x"78ffc348",
   136 => x"1ec04bd3",
   137 => x"c1f0ffc0",
   138 => x"ccfc49c1",
   139 => x"7086c487",
   140 => x"87ca0598",
   141 => x"c348d4ff",
   142 => x"48c178ff",
   143 => x"f1fd87cb",
   144 => x"058bc187",
   145 => x"c087dbff",
   146 => x"87e9fb48",
   147 => x"5c5b5e0e",
   148 => x"4cd4ff0e",
   149 => x"c687dbfd",
   150 => x"e1c01eea",
   151 => x"49c8c1f0",
   152 => x"c487d6fb",
   153 => x"02a8c186",
   154 => x"eafe87c8",
   155 => x"c148c087",
   156 => x"d2fa87e2",
   157 => x"cf497087",
   158 => x"c699ffff",
   159 => x"c802a9ea",
   160 => x"87d3fe87",
   161 => x"cbc148c0",
   162 => x"7cffc387",
   163 => x"fc4bf1c0",
   164 => x"987087f4",
   165 => x"87ebc002",
   166 => x"ffc01ec0",
   167 => x"49fac1f0",
   168 => x"c487d6fa",
   169 => x"05987086",
   170 => x"ffc387d9",
   171 => x"c3496c7c",
   172 => x"7c7c7cff",
   173 => x"99c0c17c",
   174 => x"c187c402",
   175 => x"c087d548",
   176 => x"c287d148",
   177 => x"87c405ab",
   178 => x"87c848c0",
   179 => x"fe058bc1",
   180 => x"48c087fd",
   181 => x"1e87dcf9",
   182 => x"dac21e73",
   183 => x"78c148d8",
   184 => x"d0ff4bc7",
   185 => x"fb78c248",
   186 => x"d0ff87c8",
   187 => x"c078c348",
   188 => x"d0e5c01e",
   189 => x"f849c0c1",
   190 => x"86c487ff",
   191 => x"c105a8c1",
   192 => x"abc24b87",
   193 => x"c087c505",
   194 => x"87f9c048",
   195 => x"ff058bc1",
   196 => x"f7fc87d0",
   197 => x"dcdac287",
   198 => x"05987058",
   199 => x"1ec187cd",
   200 => x"c1f0ffc0",
   201 => x"d0f849d0",
   202 => x"ff86c487",
   203 => x"ffc348d4",
   204 => x"87ddc478",
   205 => x"58e0dac2",
   206 => x"c248d0ff",
   207 => x"48d4ff78",
   208 => x"c178ffc3",
   209 => x"87edf748",
   210 => x"5c5b5e0e",
   211 => x"4a710e5d",
   212 => x"ff4dffc3",
   213 => x"7c754cd4",
   214 => x"c448d0ff",
   215 => x"7c7578c3",
   216 => x"ffc01e72",
   217 => x"49d8c1f0",
   218 => x"c487cef7",
   219 => x"02987086",
   220 => x"48c187c5",
   221 => x"7587eec0",
   222 => x"7cfec37c",
   223 => x"d41ec0c8",
   224 => x"f2f44966",
   225 => x"7586c487",
   226 => x"757c757c",
   227 => x"e0dad87c",
   228 => x"6c7c754b",
   229 => x"c187c505",
   230 => x"87f5058b",
   231 => x"d0ff7c75",
   232 => x"c078c248",
   233 => x"87c9f648",
   234 => x"5c5b5e0e",
   235 => x"4b710e5d",
   236 => x"eec54cc0",
   237 => x"ff4adfcd",
   238 => x"ffc348d4",
   239 => x"c3486878",
   240 => x"c005a8fe",
   241 => x"d4ff87fe",
   242 => x"029b734d",
   243 => x"66d087cc",
   244 => x"f449731e",
   245 => x"86c487c8",
   246 => x"d0ff87d6",
   247 => x"78d1c448",
   248 => x"d07dffc3",
   249 => x"88c14866",
   250 => x"7058a6d4",
   251 => x"87f00598",
   252 => x"c348d4ff",
   253 => x"737878ff",
   254 => x"87c5059b",
   255 => x"d048d0ff",
   256 => x"4c4ac178",
   257 => x"fe058ac1",
   258 => x"487487ed",
   259 => x"1e87e2f4",
   260 => x"4a711e73",
   261 => x"d4ff4bc0",
   262 => x"78ffc348",
   263 => x"c448d0ff",
   264 => x"d4ff78c3",
   265 => x"78ffc348",
   266 => x"ffc01e72",
   267 => x"49d1c1f0",
   268 => x"c487c6f4",
   269 => x"05987086",
   270 => x"c0c887d2",
   271 => x"4966cc1e",
   272 => x"c487e5fd",
   273 => x"ff4b7086",
   274 => x"78c248d0",
   275 => x"e4f34873",
   276 => x"5b5e0e87",
   277 => x"c00e5d5c",
   278 => x"f0ffc01e",
   279 => x"f349c9c1",
   280 => x"1ed287d7",
   281 => x"49e0dac2",
   282 => x"c887fdfc",
   283 => x"c14cc086",
   284 => x"acb7d284",
   285 => x"c287f804",
   286 => x"bf97e0da",
   287 => x"99c0c349",
   288 => x"05a9c0c1",
   289 => x"c287e7c0",
   290 => x"bf97e7da",
   291 => x"c231d049",
   292 => x"bf97e8da",
   293 => x"7232c84a",
   294 => x"e9dac2b1",
   295 => x"b14abf97",
   296 => x"ffcf4c71",
   297 => x"c19cffff",
   298 => x"c134ca84",
   299 => x"dac287e7",
   300 => x"49bf97e9",
   301 => x"99c631c1",
   302 => x"97eadac2",
   303 => x"b7c74abf",
   304 => x"c2b1722a",
   305 => x"bf97e5da",
   306 => x"9dcf4d4a",
   307 => x"97e6dac2",
   308 => x"9ac34abf",
   309 => x"dac232ca",
   310 => x"4bbf97e7",
   311 => x"b27333c2",
   312 => x"97e8dac2",
   313 => x"c0c34bbf",
   314 => x"2bb7c69b",
   315 => x"81c2b273",
   316 => x"307148c1",
   317 => x"48c14970",
   318 => x"4d703075",
   319 => x"84c14c72",
   320 => x"c0c89471",
   321 => x"cc06adb7",
   322 => x"b734c187",
   323 => x"b7c0c82d",
   324 => x"f4ff01ad",
   325 => x"f0487487",
   326 => x"5e0e87d7",
   327 => x"0e5d5c5b",
   328 => x"e3c286f8",
   329 => x"78c048c6",
   330 => x"1efedac2",
   331 => x"defb49c0",
   332 => x"7086c487",
   333 => x"87c50598",
   334 => x"c0c948c0",
   335 => x"c14dc087",
   336 => x"ddf2c07e",
   337 => x"dbc249bf",
   338 => x"c8714af4",
   339 => x"87d9ec4b",
   340 => x"c2059870",
   341 => x"c07ec087",
   342 => x"49bfd9f2",
   343 => x"4ad0dcc2",
   344 => x"ec4bc871",
   345 => x"987087c3",
   346 => x"c087c205",
   347 => x"c0026e7e",
   348 => x"e2c287fd",
   349 => x"c24dbfc4",
   350 => x"bf9ffce2",
   351 => x"d6c5487e",
   352 => x"c705a8ea",
   353 => x"c4e2c287",
   354 => x"87ce4dbf",
   355 => x"e9ca486e",
   356 => x"c502a8d5",
   357 => x"c748c087",
   358 => x"dac287e3",
   359 => x"49751efe",
   360 => x"c487ecf9",
   361 => x"05987086",
   362 => x"48c087c5",
   363 => x"c087cec7",
   364 => x"49bfd9f2",
   365 => x"4ad0dcc2",
   366 => x"ea4bc871",
   367 => x"987087eb",
   368 => x"c287c805",
   369 => x"c148c6e3",
   370 => x"c087da78",
   371 => x"49bfddf2",
   372 => x"4af4dbc2",
   373 => x"ea4bc871",
   374 => x"987087cf",
   375 => x"87c5c002",
   376 => x"d8c648c0",
   377 => x"fce2c287",
   378 => x"c149bf97",
   379 => x"c005a9d5",
   380 => x"e2c287cd",
   381 => x"49bf97fd",
   382 => x"02a9eac2",
   383 => x"c087c5c0",
   384 => x"87f9c548",
   385 => x"97fedac2",
   386 => x"c3487ebf",
   387 => x"c002a8e9",
   388 => x"486e87ce",
   389 => x"02a8ebc3",
   390 => x"c087c5c0",
   391 => x"87ddc548",
   392 => x"97c9dbc2",
   393 => x"059949bf",
   394 => x"c287ccc0",
   395 => x"bf97cadb",
   396 => x"02a9c249",
   397 => x"c087c5c0",
   398 => x"87c1c548",
   399 => x"97cbdbc2",
   400 => x"e3c248bf",
   401 => x"4c7058c2",
   402 => x"c288c148",
   403 => x"c258c6e3",
   404 => x"bf97ccdb",
   405 => x"c2817549",
   406 => x"bf97cddb",
   407 => x"7232c84a",
   408 => x"e7c27ea1",
   409 => x"786e48d3",
   410 => x"97cedbc2",
   411 => x"a6c848bf",
   412 => x"c6e3c258",
   413 => x"cfc202bf",
   414 => x"d9f2c087",
   415 => x"dcc249bf",
   416 => x"c8714ad0",
   417 => x"87e1e74b",
   418 => x"c0029870",
   419 => x"48c087c5",
   420 => x"c287eac3",
   421 => x"4cbffee2",
   422 => x"5ce7e7c2",
   423 => x"97e3dbc2",
   424 => x"31c849bf",
   425 => x"97e2dbc2",
   426 => x"49a14abf",
   427 => x"97e4dbc2",
   428 => x"32d04abf",
   429 => x"c249a172",
   430 => x"bf97e5db",
   431 => x"7232d84a",
   432 => x"66c449a1",
   433 => x"d3e7c291",
   434 => x"e7c281bf",
   435 => x"dbc259db",
   436 => x"4abf97eb",
   437 => x"dbc232c8",
   438 => x"4bbf97ea",
   439 => x"dbc24aa2",
   440 => x"4bbf97ec",
   441 => x"a27333d0",
   442 => x"eddbc24a",
   443 => x"cf4bbf97",
   444 => x"7333d89b",
   445 => x"e7c24aa2",
   446 => x"8ac25adf",
   447 => x"e7c29274",
   448 => x"a17248df",
   449 => x"87c1c178",
   450 => x"97d0dbc2",
   451 => x"31c849bf",
   452 => x"97cfdbc2",
   453 => x"49a14abf",
   454 => x"ffc731c5",
   455 => x"c229c981",
   456 => x"c259e7e7",
   457 => x"bf97d5db",
   458 => x"c232c84a",
   459 => x"bf97d4db",
   460 => x"c44aa24b",
   461 => x"826e9266",
   462 => x"5ae3e7c2",
   463 => x"48dbe7c2",
   464 => x"e7c278c0",
   465 => x"a17248d7",
   466 => x"e7e7c278",
   467 => x"dbe7c248",
   468 => x"e7c278bf",
   469 => x"e7c248eb",
   470 => x"c278bfdf",
   471 => x"02bfc6e3",
   472 => x"7487c9c0",
   473 => x"7030c448",
   474 => x"87c9c07e",
   475 => x"bfe3e7c2",
   476 => x"7030c448",
   477 => x"cae3c27e",
   478 => x"c1786e48",
   479 => x"268ef848",
   480 => x"264c264d",
   481 => x"0e4f264b",
   482 => x"5d5c5b5e",
   483 => x"c24a710e",
   484 => x"02bfc6e3",
   485 => x"4b7287cb",
   486 => x"4d722bc7",
   487 => x"c99dffc1",
   488 => x"c84b7287",
   489 => x"c34d722b",
   490 => x"e7c29dff",
   491 => x"c083bfd3",
   492 => x"abbfd5f2",
   493 => x"c087d902",
   494 => x"c25bd9f2",
   495 => x"731efeda",
   496 => x"87cbf149",
   497 => x"987086c4",
   498 => x"c087c505",
   499 => x"87e6c048",
   500 => x"bfc6e3c2",
   501 => x"7587d202",
   502 => x"c291c449",
   503 => x"6981feda",
   504 => x"ffffcf4c",
   505 => x"cb9cffff",
   506 => x"c2497587",
   507 => x"fedac291",
   508 => x"4c699f81",
   509 => x"c6fe4874",
   510 => x"5b5e0e87",
   511 => x"f80e5d5c",
   512 => x"9c4c7186",
   513 => x"c087c505",
   514 => x"87c0c348",
   515 => x"487ea4c8",
   516 => x"66d878c0",
   517 => x"d887c702",
   518 => x"05bf9766",
   519 => x"48c087c5",
   520 => x"c087e9c2",
   521 => x"4949c11e",
   522 => x"c487d3ca",
   523 => x"9d4d7086",
   524 => x"87c2c102",
   525 => x"4acee3c2",
   526 => x"e04966d8",
   527 => x"987087d0",
   528 => x"87f2c002",
   529 => x"66d84a75",
   530 => x"e04bcb49",
   531 => x"987087f5",
   532 => x"87e2c002",
   533 => x"9d751ec0",
   534 => x"c887c702",
   535 => x"78c048a6",
   536 => x"a6c887c5",
   537 => x"c878c148",
   538 => x"d1c94966",
   539 => x"7086c487",
   540 => x"fe059d4d",
   541 => x"9d7587fe",
   542 => x"87cec102",
   543 => x"6e49a5dc",
   544 => x"da786948",
   545 => x"a6c449a5",
   546 => x"78a4c448",
   547 => x"c448699f",
   548 => x"c2780866",
   549 => x"02bfc6e3",
   550 => x"a5d487d2",
   551 => x"49699f49",
   552 => x"99ffffc0",
   553 => x"30d04871",
   554 => x"87c27e70",
   555 => x"486e7ec0",
   556 => x"80bf66c4",
   557 => x"780866c4",
   558 => x"a4cc7cc0",
   559 => x"bf66c449",
   560 => x"49a4d079",
   561 => x"48c179c0",
   562 => x"48c087c2",
   563 => x"eefa8ef8",
   564 => x"5b5e0e87",
   565 => x"4c710e5c",
   566 => x"cbc1029c",
   567 => x"49a4c887",
   568 => x"c3c10269",
   569 => x"cc496c87",
   570 => x"80714866",
   571 => x"7058a6d0",
   572 => x"c2e3c2b9",
   573 => x"baff4abf",
   574 => x"99719972",
   575 => x"87e5c002",
   576 => x"6b4ba4c4",
   577 => x"87fff949",
   578 => x"e2c27b70",
   579 => x"6c49bffe",
   580 => x"cc7c7181",
   581 => x"e3c2b966",
   582 => x"ff4abfc2",
   583 => x"719972ba",
   584 => x"dbff0599",
   585 => x"7c66cc87",
   586 => x"1e87d6f9",
   587 => x"4b711e73",
   588 => x"87c7029b",
   589 => x"6949a3c8",
   590 => x"c087c505",
   591 => x"87f6c048",
   592 => x"bfd7e7c2",
   593 => x"4aa3c449",
   594 => x"8ac24a6a",
   595 => x"bffee2c2",
   596 => x"49a17292",
   597 => x"bfc2e3c2",
   598 => x"729a6b4a",
   599 => x"f2c049a1",
   600 => x"66c859d9",
   601 => x"e6ea711e",
   602 => x"7086c487",
   603 => x"87c40598",
   604 => x"87c248c0",
   605 => x"caf848c1",
   606 => x"1e731e87",
   607 => x"029b4b71",
   608 => x"a3c887c7",
   609 => x"c5056949",
   610 => x"c048c087",
   611 => x"e7c287f6",
   612 => x"c449bfd7",
   613 => x"4a6a4aa3",
   614 => x"e2c28ac2",
   615 => x"7292bffe",
   616 => x"e3c249a1",
   617 => x"6b4abfc2",
   618 => x"49a1729a",
   619 => x"59d9f2c0",
   620 => x"711e66c8",
   621 => x"c487d1e6",
   622 => x"05987086",
   623 => x"48c087c4",
   624 => x"48c187c2",
   625 => x"0e87fcf6",
   626 => x"5d5c5b5e",
   627 => x"4b711e0e",
   628 => x"734d66d4",
   629 => x"ccc1029b",
   630 => x"49a3c887",
   631 => x"c4c10269",
   632 => x"4ca3d087",
   633 => x"bfc2e3c2",
   634 => x"6cb9ff49",
   635 => x"d47e994a",
   636 => x"cd06a966",
   637 => x"7c7bc087",
   638 => x"c44aa3cc",
   639 => x"796a49a3",
   640 => x"497287ca",
   641 => x"d499c0f8",
   642 => x"8d714d66",
   643 => x"29c94975",
   644 => x"49731e71",
   645 => x"c287fafa",
   646 => x"731efeda",
   647 => x"87cbfc49",
   648 => x"66d486c8",
   649 => x"d6f5267c",
   650 => x"1e731e87",
   651 => x"029b4b71",
   652 => x"c287e4c0",
   653 => x"735bebe7",
   654 => x"c28ac24a",
   655 => x"49bffee2",
   656 => x"d7e7c292",
   657 => x"807248bf",
   658 => x"58efe7c2",
   659 => x"30c44871",
   660 => x"58cee3c2",
   661 => x"c287edc0",
   662 => x"c248e7e7",
   663 => x"78bfdbe7",
   664 => x"48ebe7c2",
   665 => x"bfdfe7c2",
   666 => x"c6e3c278",
   667 => x"87c902bf",
   668 => x"bffee2c2",
   669 => x"c731c449",
   670 => x"e3e7c287",
   671 => x"31c449bf",
   672 => x"59cee3c2",
   673 => x"0e87fcf3",
   674 => x"0e5c5b5e",
   675 => x"4bc04a71",
   676 => x"c0029a72",
   677 => x"a2da87e0",
   678 => x"4b699f49",
   679 => x"bfc6e3c2",
   680 => x"d487cf02",
   681 => x"699f49a2",
   682 => x"ffc04c49",
   683 => x"34d09cff",
   684 => x"4cc087c2",
   685 => x"4973b374",
   686 => x"f387eefd",
   687 => x"5e0e87c3",
   688 => x"0e5d5c5b",
   689 => x"4a7186f4",
   690 => x"9a727ec0",
   691 => x"c287d802",
   692 => x"c048fada",
   693 => x"f2dac278",
   694 => x"ebe7c248",
   695 => x"dac278bf",
   696 => x"e7c248f6",
   697 => x"c278bfe7",
   698 => x"c048dbe3",
   699 => x"cae3c250",
   700 => x"dac249bf",
   701 => x"714abffa",
   702 => x"c9c403aa",
   703 => x"cf497287",
   704 => x"e9c00599",
   705 => x"d5f2c087",
   706 => x"f2dac248",
   707 => x"dac278bf",
   708 => x"dac21efe",
   709 => x"c249bff2",
   710 => x"c148f2da",
   711 => x"e37178a1",
   712 => x"86c487ed",
   713 => x"48d1f2c0",
   714 => x"78fedac2",
   715 => x"f2c087cc",
   716 => x"c048bfd1",
   717 => x"f2c080e0",
   718 => x"dac258d5",
   719 => x"c148bffa",
   720 => x"fedac280",
   721 => x"0c912758",
   722 => x"97bf0000",
   723 => x"029d4dbf",
   724 => x"c387e3c2",
   725 => x"c202ade5",
   726 => x"f2c087dc",
   727 => x"cb4bbfd1",
   728 => x"4c1149a3",
   729 => x"c105accf",
   730 => x"497587d2",
   731 => x"89c199df",
   732 => x"e3c291cd",
   733 => x"a3c181ce",
   734 => x"c351124a",
   735 => x"51124aa3",
   736 => x"124aa3c5",
   737 => x"4aa3c751",
   738 => x"a3c95112",
   739 => x"ce51124a",
   740 => x"51124aa3",
   741 => x"124aa3d0",
   742 => x"4aa3d251",
   743 => x"a3d45112",
   744 => x"d651124a",
   745 => x"51124aa3",
   746 => x"124aa3d8",
   747 => x"4aa3dc51",
   748 => x"a3de5112",
   749 => x"c151124a",
   750 => x"87fac07e",
   751 => x"99c84974",
   752 => x"87ebc005",
   753 => x"99d04974",
   754 => x"dc87d105",
   755 => x"cbc00266",
   756 => x"dc497387",
   757 => x"98700f66",
   758 => x"87d3c002",
   759 => x"c6c0056e",
   760 => x"cee3c287",
   761 => x"c050c048",
   762 => x"48bfd1f2",
   763 => x"c287ddc2",
   764 => x"c048dbe3",
   765 => x"e3c27e50",
   766 => x"c249bfca",
   767 => x"4abffada",
   768 => x"fb04aa71",
   769 => x"e7c287f7",
   770 => x"c005bfeb",
   771 => x"e3c287c8",
   772 => x"c102bfc6",
   773 => x"dac287f4",
   774 => x"ed49bff6",
   775 => x"dac287e9",
   776 => x"a6c458fa",
   777 => x"f6dac248",
   778 => x"e3c278bf",
   779 => x"c002bfc6",
   780 => x"66c487d8",
   781 => x"ffffcf49",
   782 => x"a999f8ff",
   783 => x"87c5c002",
   784 => x"e1c04cc0",
   785 => x"c04cc187",
   786 => x"66c487dc",
   787 => x"f8ffcf49",
   788 => x"c002a999",
   789 => x"a6c887c8",
   790 => x"c078c048",
   791 => x"a6c887c5",
   792 => x"c878c148",
   793 => x"9c744c66",
   794 => x"87dec005",
   795 => x"c24966c4",
   796 => x"fee2c289",
   797 => x"e7c291bf",
   798 => x"7148bfd7",
   799 => x"f6dac280",
   800 => x"fadac258",
   801 => x"f978c048",
   802 => x"48c087e3",
   803 => x"eeeb8ef4",
   804 => x"00000087",
   805 => x"ffffff00",
   806 => x"000ca1ff",
   807 => x"000caa00",
   808 => x"54414600",
   809 => x"20203233",
   810 => x"41460020",
   811 => x"20363154",
   812 => x"1e002020",
   813 => x"c348d4ff",
   814 => x"486878ff",
   815 => x"ff1e4f26",
   816 => x"ffc348d4",
   817 => x"48d0ff78",
   818 => x"ff78e1c0",
   819 => x"78d448d4",
   820 => x"48efe7c2",
   821 => x"50bfd4ff",
   822 => x"ff1e4f26",
   823 => x"e0c048d0",
   824 => x"1e4f2678",
   825 => x"7087ccff",
   826 => x"c6029949",
   827 => x"a9fbc087",
   828 => x"7187f105",
   829 => x"0e4f2648",
   830 => x"0e5c5b5e",
   831 => x"4cc04b71",
   832 => x"7087f0fe",
   833 => x"c0029949",
   834 => x"ecc087f9",
   835 => x"f2c002a9",
   836 => x"a9fbc087",
   837 => x"87ebc002",
   838 => x"acb766cc",
   839 => x"d087c703",
   840 => x"87c20266",
   841 => x"99715371",
   842 => x"c187c202",
   843 => x"87c3fe84",
   844 => x"02994970",
   845 => x"ecc087cd",
   846 => x"87c702a9",
   847 => x"05a9fbc0",
   848 => x"d087d5ff",
   849 => x"87c30266",
   850 => x"c07b97c0",
   851 => x"c405a9ec",
   852 => x"c54a7487",
   853 => x"c04a7487",
   854 => x"48728a0a",
   855 => x"4d2687c2",
   856 => x"4b264c26",
   857 => x"fd1e4f26",
   858 => x"4a7087c9",
   859 => x"04aaf0c0",
   860 => x"f9c087c9",
   861 => x"87c301aa",
   862 => x"c18af0c0",
   863 => x"c904aac1",
   864 => x"aadac187",
   865 => x"c087c301",
   866 => x"48728af7",
   867 => x"5e0e4f26",
   868 => x"710e5c5b",
   869 => x"4bd4ff4a",
   870 => x"e7c04972",
   871 => x"9c4c7087",
   872 => x"c187c202",
   873 => x"48d0ff8c",
   874 => x"d5c178c5",
   875 => x"c649747b",
   876 => x"eee3c131",
   877 => x"484abf97",
   878 => x"7b70b071",
   879 => x"c448d0ff",
   880 => x"87dcfe78",
   881 => x"5c5b5e0e",
   882 => x"86f80e5d",
   883 => x"7ec04c71",
   884 => x"c087ebfb",
   885 => x"f1f9c04b",
   886 => x"c049bf97",
   887 => x"87cf04a9",
   888 => x"c187c0fc",
   889 => x"f1f9c083",
   890 => x"ab49bf97",
   891 => x"c087f106",
   892 => x"bf97f1f9",
   893 => x"fa87cf02",
   894 => x"497087f9",
   895 => x"87c60299",
   896 => x"05a9ecc0",
   897 => x"4bc087f1",
   898 => x"7087e8fa",
   899 => x"87e3fa4d",
   900 => x"fa58a6c8",
   901 => x"4a7087dd",
   902 => x"a4c883c1",
   903 => x"49699749",
   904 => x"87c702ad",
   905 => x"05adffc0",
   906 => x"c987e7c0",
   907 => x"699749a4",
   908 => x"a966c449",
   909 => x"4887c702",
   910 => x"05a8ffc0",
   911 => x"a4ca87d4",
   912 => x"49699749",
   913 => x"87c602aa",
   914 => x"05aaffc0",
   915 => x"7ec187c4",
   916 => x"ecc087d0",
   917 => x"87c602ad",
   918 => x"05adfbc0",
   919 => x"4bc087c4",
   920 => x"026e7ec1",
   921 => x"f987e1fe",
   922 => x"487387f0",
   923 => x"edfb8ef8",
   924 => x"5e0e0087",
   925 => x"0e5d5c5b",
   926 => x"4d7186f8",
   927 => x"754bd4ff",
   928 => x"f4e7c21e",
   929 => x"87f1e549",
   930 => x"987086c4",
   931 => x"87cac402",
   932 => x"c148a6c4",
   933 => x"78bff0e3",
   934 => x"f1fb4975",
   935 => x"48d0ff87",
   936 => x"d6c178c5",
   937 => x"754ac07b",
   938 => x"7b1149a2",
   939 => x"b7cb82c1",
   940 => x"87f304aa",
   941 => x"ffc34acc",
   942 => x"c082c17b",
   943 => x"04aab7e0",
   944 => x"d0ff87f4",
   945 => x"c378c448",
   946 => x"78c57bff",
   947 => x"c17bd3c1",
   948 => x"6678c47b",
   949 => x"a8b7c048",
   950 => x"87eec206",
   951 => x"bffce7c2",
   952 => x"4866c44c",
   953 => x"a6c88874",
   954 => x"029c7458",
   955 => x"c287f7c1",
   956 => x"c87efeda",
   957 => x"c08c4dc0",
   958 => x"c603acb7",
   959 => x"a4c0c887",
   960 => x"c24cc04d",
   961 => x"bf97efe7",
   962 => x"0299d049",
   963 => x"1ec087d0",
   964 => x"49f4e7c2",
   965 => x"c487d4e8",
   966 => x"c04a7086",
   967 => x"dac287ed",
   968 => x"e7c21efe",
   969 => x"c2e849f4",
   970 => x"7086c487",
   971 => x"48d0ff4a",
   972 => x"c178c5c8",
   973 => x"976e7bd4",
   974 => x"486e7bbf",
   975 => x"7e7080c1",
   976 => x"ff058dc1",
   977 => x"d0ff87f0",
   978 => x"7278c448",
   979 => x"87c5059a",
   980 => x"c7c148c0",
   981 => x"c21ec187",
   982 => x"e549f4e7",
   983 => x"86c487f3",
   984 => x"fe059c74",
   985 => x"66c487c9",
   986 => x"a8b7c048",
   987 => x"c287d106",
   988 => x"c048f4e7",
   989 => x"c080d078",
   990 => x"c280f478",
   991 => x"78bfc0e8",
   992 => x"c04866c4",
   993 => x"fd01a8b7",
   994 => x"d0ff87d2",
   995 => x"c178c548",
   996 => x"7bc07bd3",
   997 => x"48c178c4",
   998 => x"48c087c2",
   999 => x"4d268ef8",
  1000 => x"4b264c26",
  1001 => x"5e0e4f26",
  1002 => x"0e5d5c5b",
  1003 => x"c04b711e",
  1004 => x"04ab4d4c",
  1005 => x"c087e8c0",
  1006 => x"751ec4f7",
  1007 => x"87c4029d",
  1008 => x"87c24ac0",
  1009 => x"49724ac1",
  1010 => x"c487f3eb",
  1011 => x"c17e7086",
  1012 => x"c2056e84",
  1013 => x"c14c7387",
  1014 => x"06ac7385",
  1015 => x"6e87d8ff",
  1016 => x"f9fe2648",
  1017 => x"5b5e0e87",
  1018 => x"4b710e5c",
  1019 => x"d80266cc",
  1020 => x"f0c04c87",
  1021 => x"87d8028c",
  1022 => x"8ac14a74",
  1023 => x"8a87d102",
  1024 => x"8a87cd02",
  1025 => x"d987c902",
  1026 => x"f9497387",
  1027 => x"87d287e4",
  1028 => x"49c01e74",
  1029 => x"87f5d7c1",
  1030 => x"49731e74",
  1031 => x"87edd7c1",
  1032 => x"fbfd86c8",
  1033 => x"5b5e0e87",
  1034 => x"1e0e5d5c",
  1035 => x"de494c71",
  1036 => x"dce8c291",
  1037 => x"9785714d",
  1038 => x"dcc1026d",
  1039 => x"c8e8c287",
  1040 => x"817449bf",
  1041 => x"87defd71",
  1042 => x"98487e70",
  1043 => x"87f2c002",
  1044 => x"4bd0e8c2",
  1045 => x"49cb4a70",
  1046 => x"87cbc1ff",
  1047 => x"93cb4b74",
  1048 => x"83c2e4c1",
  1049 => x"c2c183c4",
  1050 => x"49747bdd",
  1051 => x"87cbc1c1",
  1052 => x"e3c17b75",
  1053 => x"49bf97ef",
  1054 => x"d0e8c21e",
  1055 => x"87e5fd49",
  1056 => x"497486c4",
  1057 => x"87f3c0c1",
  1058 => x"c2c149c0",
  1059 => x"e7c287d2",
  1060 => x"78c048f0",
  1061 => x"fbdd49c1",
  1062 => x"c1fc2687",
  1063 => x"616f4c87",
  1064 => x"676e6964",
  1065 => x"002e2e2e",
  1066 => x"711e731e",
  1067 => x"e8c2494a",
  1068 => x"7181bfc8",
  1069 => x"7087effb",
  1070 => x"c4029b4b",
  1071 => x"c6e74987",
  1072 => x"c8e8c287",
  1073 => x"c178c048",
  1074 => x"87c8dd49",
  1075 => x"1e87d3fb",
  1076 => x"c1c149c0",
  1077 => x"4f2687ca",
  1078 => x"494a711e",
  1079 => x"e4c191cb",
  1080 => x"81c881c2",
  1081 => x"e7c24811",
  1082 => x"e8c258f4",
  1083 => x"78c048c8",
  1084 => x"dfdc49c1",
  1085 => x"1e4f2687",
  1086 => x"d2029971",
  1087 => x"d7e5c187",
  1088 => x"f750c048",
  1089 => x"d8c3c180",
  1090 => x"fbe3c140",
  1091 => x"c187ce78",
  1092 => x"c148d3e5",
  1093 => x"fc78f4e3",
  1094 => x"cfc3c180",
  1095 => x"0e4f2678",
  1096 => x"5d5c5b5e",
  1097 => x"c286f40e",
  1098 => x"c04dfeda",
  1099 => x"48a6c44c",
  1100 => x"e8c278c0",
  1101 => x"c048bfc8",
  1102 => x"c0c106a8",
  1103 => x"fedac287",
  1104 => x"c0029848",
  1105 => x"f7c087f7",
  1106 => x"66c81ec4",
  1107 => x"c487c702",
  1108 => x"78c048a6",
  1109 => x"a6c487c5",
  1110 => x"c478c148",
  1111 => x"dde54966",
  1112 => x"7086c487",
  1113 => x"c484c14d",
  1114 => x"80c14866",
  1115 => x"c258a6c8",
  1116 => x"acbfc8e8",
  1117 => x"7587c603",
  1118 => x"c9ff059d",
  1119 => x"754cc087",
  1120 => x"dcc3029d",
  1121 => x"c4f7c087",
  1122 => x"0266c81e",
  1123 => x"a6cc87c7",
  1124 => x"c578c048",
  1125 => x"48a6cc87",
  1126 => x"66cc78c1",
  1127 => x"87dee449",
  1128 => x"7e7086c4",
  1129 => x"c2029848",
  1130 => x"cb4987e4",
  1131 => x"49699781",
  1132 => x"c10299d0",
  1133 => x"497487d4",
  1134 => x"e4c191cb",
  1135 => x"c2c181c2",
  1136 => x"81c879e8",
  1137 => x"7451ffc3",
  1138 => x"c291de49",
  1139 => x"714ddce8",
  1140 => x"97c1c285",
  1141 => x"49a5c17d",
  1142 => x"c251e0c0",
  1143 => x"bf97cee3",
  1144 => x"c187d202",
  1145 => x"4ba5c284",
  1146 => x"4acee3c2",
  1147 => x"fafe49db",
  1148 => x"d9c187f5",
  1149 => x"49a5cd87",
  1150 => x"84c151c0",
  1151 => x"6e4ba5c2",
  1152 => x"fe49cb4a",
  1153 => x"c187e0fa",
  1154 => x"497487c4",
  1155 => x"e4c191cb",
  1156 => x"c0c181c2",
  1157 => x"e3c279e5",
  1158 => x"02bf97ce",
  1159 => x"497487d8",
  1160 => x"84c191de",
  1161 => x"4bdce8c2",
  1162 => x"e3c28371",
  1163 => x"49dd4ace",
  1164 => x"87f3f9fe",
  1165 => x"4b7487d8",
  1166 => x"e8c293de",
  1167 => x"a3cb83dc",
  1168 => x"c151c049",
  1169 => x"4a6e7384",
  1170 => x"f9fe49cb",
  1171 => x"66c487d9",
  1172 => x"c880c148",
  1173 => x"acc758a6",
  1174 => x"87c5c003",
  1175 => x"e4fc056e",
  1176 => x"f4487487",
  1177 => x"87f6f48e",
  1178 => x"711e731e",
  1179 => x"91cb494b",
  1180 => x"81c2e4c1",
  1181 => x"c14aa1c8",
  1182 => x"1248eee3",
  1183 => x"4aa1c950",
  1184 => x"48f1f9c0",
  1185 => x"81ca5012",
  1186 => x"48efe3c1",
  1187 => x"e3c15011",
  1188 => x"49bf97ef",
  1189 => x"f549c01e",
  1190 => x"e7c287cb",
  1191 => x"78de48f0",
  1192 => x"efd549c1",
  1193 => x"f9f32687",
  1194 => x"5b5e0e87",
  1195 => x"f40e5d5c",
  1196 => x"494d7186",
  1197 => x"e4c191cb",
  1198 => x"a1c881c2",
  1199 => x"7ea1ca4a",
  1200 => x"c248a6c4",
  1201 => x"78bff8eb",
  1202 => x"4bbf976e",
  1203 => x"734c66c4",
  1204 => x"cc48122c",
  1205 => x"9c7058a6",
  1206 => x"81c984c1",
  1207 => x"b7496997",
  1208 => x"87c204ac",
  1209 => x"976e4cc0",
  1210 => x"66c84abf",
  1211 => x"ff317249",
  1212 => x"9966c4b9",
  1213 => x"30724874",
  1214 => x"71484a70",
  1215 => x"fcebc2b0",
  1216 => x"f6e4c058",
  1217 => x"d449c087",
  1218 => x"497587ca",
  1219 => x"87ebf6c0",
  1220 => x"c9f28ef4",
  1221 => x"1e731e87",
  1222 => x"fe494b71",
  1223 => x"497387cb",
  1224 => x"f187c6fe",
  1225 => x"731e87fc",
  1226 => x"c64b711e",
  1227 => x"db024aa3",
  1228 => x"028ac187",
  1229 => x"028a87d6",
  1230 => x"8a87dac1",
  1231 => x"87fcc002",
  1232 => x"e1c0028a",
  1233 => x"cb028a87",
  1234 => x"87dbc187",
  1235 => x"c7f649c7",
  1236 => x"87dec187",
  1237 => x"bfc8e8c2",
  1238 => x"87cbc102",
  1239 => x"c288c148",
  1240 => x"c158cce8",
  1241 => x"e8c287c1",
  1242 => x"c002bfcc",
  1243 => x"e8c287f9",
  1244 => x"c148bfc8",
  1245 => x"cce8c280",
  1246 => x"87ebc058",
  1247 => x"bfc8e8c2",
  1248 => x"c289c649",
  1249 => x"c059cce8",
  1250 => x"da03a9b7",
  1251 => x"c8e8c287",
  1252 => x"d278c048",
  1253 => x"cce8c287",
  1254 => x"87cb02bf",
  1255 => x"bfc8e8c2",
  1256 => x"c280c648",
  1257 => x"c058cce8",
  1258 => x"87e8d149",
  1259 => x"f4c04973",
  1260 => x"edef87c9",
  1261 => x"5b5e0e87",
  1262 => x"ff0e5d5c",
  1263 => x"a6dc86d4",
  1264 => x"48a6c859",
  1265 => x"80c478c0",
  1266 => x"7866c0c1",
  1267 => x"78c180c4",
  1268 => x"78c180c4",
  1269 => x"48cce8c2",
  1270 => x"e7c278c1",
  1271 => x"de48bff0",
  1272 => x"87c905a8",
  1273 => x"cc87f8f4",
  1274 => x"e6cf58a6",
  1275 => x"87cee387",
  1276 => x"e287f0e3",
  1277 => x"4c7087fd",
  1278 => x"02acfbc0",
  1279 => x"d887fbc1",
  1280 => x"edc10566",
  1281 => x"66fcc087",
  1282 => x"6a82c44a",
  1283 => x"c11e727e",
  1284 => x"c448c8e0",
  1285 => x"a1c84966",
  1286 => x"7141204a",
  1287 => x"87f905aa",
  1288 => x"4a265110",
  1289 => x"4866fcc0",
  1290 => x"78e8c9c1",
  1291 => x"81c7496a",
  1292 => x"fcc05174",
  1293 => x"81c84966",
  1294 => x"fcc051c1",
  1295 => x"81c94966",
  1296 => x"fcc051c0",
  1297 => x"81ca4966",
  1298 => x"1ec151c0",
  1299 => x"496a1ed8",
  1300 => x"e2e281c8",
  1301 => x"c186c887",
  1302 => x"c04866c0",
  1303 => x"87c701a8",
  1304 => x"c148a6c8",
  1305 => x"c187ce78",
  1306 => x"c14866c0",
  1307 => x"58a6d088",
  1308 => x"eee187c3",
  1309 => x"48a6d087",
  1310 => x"9c7478c2",
  1311 => x"87cfcd02",
  1312 => x"c14866c8",
  1313 => x"03a866c4",
  1314 => x"dc87c4cd",
  1315 => x"78c048a6",
  1316 => x"78c080e8",
  1317 => x"7087dce0",
  1318 => x"acd0c14c",
  1319 => x"87d7c205",
  1320 => x"e37e66c4",
  1321 => x"a6c887c0",
  1322 => x"87c7e058",
  1323 => x"ecc04c70",
  1324 => x"edc105ac",
  1325 => x"4966c887",
  1326 => x"fcc091cb",
  1327 => x"a1c48166",
  1328 => x"c84d6a4a",
  1329 => x"66c44aa1",
  1330 => x"d8c3c152",
  1331 => x"e2dfff79",
  1332 => x"9c4c7087",
  1333 => x"c087d902",
  1334 => x"d302acfb",
  1335 => x"ff557487",
  1336 => x"7087d0df",
  1337 => x"c7029c4c",
  1338 => x"acfbc087",
  1339 => x"87edff05",
  1340 => x"c255e0c0",
  1341 => x"97c055c1",
  1342 => x"4866d87d",
  1343 => x"db05a86e",
  1344 => x"4866c887",
  1345 => x"04a866cc",
  1346 => x"66c887ca",
  1347 => x"cc80c148",
  1348 => x"87c858a6",
  1349 => x"c14866cc",
  1350 => x"58a6d088",
  1351 => x"87d3deff",
  1352 => x"d0c14c70",
  1353 => x"87c805ac",
  1354 => x"c14866d4",
  1355 => x"58a6d880",
  1356 => x"02acd0c1",
  1357 => x"c487e9fd",
  1358 => x"66d84866",
  1359 => x"e0c905a8",
  1360 => x"a6e0c087",
  1361 => x"7478c048",
  1362 => x"88fbc048",
  1363 => x"98487e70",
  1364 => x"87e2c902",
  1365 => x"7088cb48",
  1366 => x"0298487e",
  1367 => x"4887cdc1",
  1368 => x"7e7088c9",
  1369 => x"c3029848",
  1370 => x"c44887fe",
  1371 => x"487e7088",
  1372 => x"87ce0298",
  1373 => x"7088c148",
  1374 => x"0298487e",
  1375 => x"c887e9c3",
  1376 => x"a6dc87d6",
  1377 => x"78f0c048",
  1378 => x"87e7dcff",
  1379 => x"ecc04c70",
  1380 => x"c4c002ac",
  1381 => x"a6e0c087",
  1382 => x"acecc05c",
  1383 => x"ff87cd02",
  1384 => x"7087d0dc",
  1385 => x"acecc04c",
  1386 => x"87f3ff05",
  1387 => x"02acecc0",
  1388 => x"ff87c4c0",
  1389 => x"c087fcdb",
  1390 => x"d01eca1e",
  1391 => x"91cb4966",
  1392 => x"4866c4c1",
  1393 => x"a6cc8071",
  1394 => x"4866c858",
  1395 => x"a6d080c4",
  1396 => x"bf66cc58",
  1397 => x"dedcff49",
  1398 => x"de1ec187",
  1399 => x"bf66d41e",
  1400 => x"d2dcff49",
  1401 => x"7086d087",
  1402 => x"08c04849",
  1403 => x"a6e8c088",
  1404 => x"06a8c058",
  1405 => x"c087eec0",
  1406 => x"dd4866e4",
  1407 => x"e4c003a8",
  1408 => x"bf66c487",
  1409 => x"66e4c049",
  1410 => x"51e0c081",
  1411 => x"4966e4c0",
  1412 => x"66c481c1",
  1413 => x"c1c281bf",
  1414 => x"66e4c051",
  1415 => x"c481c249",
  1416 => x"c081bf66",
  1417 => x"c1486e51",
  1418 => x"6e78e8c9",
  1419 => x"d081c849",
  1420 => x"496e5166",
  1421 => x"66d481c9",
  1422 => x"ca496e51",
  1423 => x"5166dc81",
  1424 => x"c14866d0",
  1425 => x"58a6d480",
  1426 => x"cc4866c8",
  1427 => x"c004a866",
  1428 => x"66c887cb",
  1429 => x"cc80c148",
  1430 => x"d9c558a6",
  1431 => x"4866cc87",
  1432 => x"a6d088c1",
  1433 => x"87cec558",
  1434 => x"87fadbff",
  1435 => x"58a6e8c0",
  1436 => x"87f2dbff",
  1437 => x"58a6e0c0",
  1438 => x"05a8ecc0",
  1439 => x"dc87cac0",
  1440 => x"e4c048a6",
  1441 => x"c4c07866",
  1442 => x"e6d8ff87",
  1443 => x"4966c887",
  1444 => x"fcc091cb",
  1445 => x"80714866",
  1446 => x"c84a7e70",
  1447 => x"ca496e82",
  1448 => x"66e4c081",
  1449 => x"4966dc51",
  1450 => x"e4c081c1",
  1451 => x"48c18966",
  1452 => x"49703071",
  1453 => x"977189c1",
  1454 => x"f8ebc27a",
  1455 => x"e4c049bf",
  1456 => x"6a972966",
  1457 => x"9871484a",
  1458 => x"58a6ecc0",
  1459 => x"81c4496e",
  1460 => x"66d84d69",
  1461 => x"a866c448",
  1462 => x"87c8c002",
  1463 => x"c048a6c4",
  1464 => x"87c5c078",
  1465 => x"c148a6c4",
  1466 => x"1e66c478",
  1467 => x"751ee0c0",
  1468 => x"c2d8ff49",
  1469 => x"7086c887",
  1470 => x"acb7c04c",
  1471 => x"87d4c106",
  1472 => x"e0c08574",
  1473 => x"75897449",
  1474 => x"d1e0c14b",
  1475 => x"e6fe714a",
  1476 => x"85c287d5",
  1477 => x"4866e0c0",
  1478 => x"e4c080c1",
  1479 => x"e8c058a6",
  1480 => x"81c14966",
  1481 => x"c002a970",
  1482 => x"a6c487c8",
  1483 => x"c078c048",
  1484 => x"a6c487c5",
  1485 => x"c478c148",
  1486 => x"a4c21e66",
  1487 => x"48e0c049",
  1488 => x"49708871",
  1489 => x"ff49751e",
  1490 => x"c887ecd6",
  1491 => x"a8b7c086",
  1492 => x"87c0ff01",
  1493 => x"0266e0c0",
  1494 => x"6e87d1c0",
  1495 => x"c081c949",
  1496 => x"6e5166e0",
  1497 => x"e9cac148",
  1498 => x"87ccc078",
  1499 => x"81c9496e",
  1500 => x"486e51c2",
  1501 => x"78d5ccc1",
  1502 => x"cc4866c8",
  1503 => x"c004a866",
  1504 => x"66c887cb",
  1505 => x"cc80c148",
  1506 => x"e9c058a6",
  1507 => x"4866cc87",
  1508 => x"a6d088c1",
  1509 => x"87dec058",
  1510 => x"87c7d5ff",
  1511 => x"d5c04c70",
  1512 => x"acc6c187",
  1513 => x"87c8c005",
  1514 => x"c14866d0",
  1515 => x"58a6d480",
  1516 => x"87efd4ff",
  1517 => x"66d44c70",
  1518 => x"d880c148",
  1519 => x"9c7458a6",
  1520 => x"87cbc002",
  1521 => x"c14866c8",
  1522 => x"04a866c4",
  1523 => x"ff87fcf2",
  1524 => x"c887c7d4",
  1525 => x"a8c74866",
  1526 => x"87e5c003",
  1527 => x"48cce8c2",
  1528 => x"66c878c0",
  1529 => x"c091cb49",
  1530 => x"c48166fc",
  1531 => x"4a6a4aa1",
  1532 => x"c87952c0",
  1533 => x"80c14866",
  1534 => x"c758a6cc",
  1535 => x"dbff04a8",
  1536 => x"8ed4ff87",
  1537 => x"87d6deff",
  1538 => x"64616f4c",
  1539 => x"202e2a20",
  1540 => x"00203a00",
  1541 => x"711e731e",
  1542 => x"c6029b4b",
  1543 => x"c8e8c287",
  1544 => x"c778c048",
  1545 => x"c8e8c21e",
  1546 => x"e4c11ebf",
  1547 => x"e7c21ec2",
  1548 => x"ed49bff0",
  1549 => x"86cc87ff",
  1550 => x"bff0e7c2",
  1551 => x"87f7e249",
  1552 => x"c8029b73",
  1553 => x"c2e4c187",
  1554 => x"c0e3c049",
  1555 => x"d1ddff87",
  1556 => x"e3c11e87",
  1557 => x"50c048ee",
  1558 => x"bfe5e5c1",
  1559 => x"d1d8ff49",
  1560 => x"2648c087",
  1561 => x"e3c71e4f",
  1562 => x"fe49c187",
  1563 => x"e9fe87e6",
  1564 => x"987087e5",
  1565 => x"fe87cd02",
  1566 => x"7087dff2",
  1567 => x"87c40298",
  1568 => x"87c24ac1",
  1569 => x"9a724ac0",
  1570 => x"c087ce05",
  1571 => x"f5e2c11e",
  1572 => x"eeeec049",
  1573 => x"fe86c487",
  1574 => x"c11ec087",
  1575 => x"c049c0e3",
  1576 => x"c087e0ee",
  1577 => x"87e9fe1e",
  1578 => x"eec04970",
  1579 => x"dac387d5",
  1580 => x"268ef887",
  1581 => x"2044534f",
  1582 => x"6c696166",
  1583 => x"002e6465",
  1584 => x"746f6f42",
  1585 => x"2e676e69",
  1586 => x"1e002e2e",
  1587 => x"87fae5c0",
  1588 => x"87e9f1c0",
  1589 => x"4f2687f6",
  1590 => x"c8e8c21e",
  1591 => x"c278c048",
  1592 => x"c048f0e7",
  1593 => x"87fdfd78",
  1594 => x"48c087e1",
  1595 => x"00004f26",
  1596 => x"00000001",
  1597 => x"78452080",
  1598 => x"80007469",
  1599 => x"63614220",
  1600 => x"1025006b",
  1601 => x"2a1c0000",
  1602 => x"00000000",
  1603 => x"00102500",
  1604 => x"002a3a00",
  1605 => x"00000000",
  1606 => x"00001025",
  1607 => x"00002a58",
  1608 => x"25000000",
  1609 => x"76000010",
  1610 => x"0000002a",
  1611 => x"10250000",
  1612 => x"2a940000",
  1613 => x"00000000",
  1614 => x"00102500",
  1615 => x"002ab200",
  1616 => x"00000000",
  1617 => x"00001025",
  1618 => x"00002ad0",
  1619 => x"d8000000",
  1620 => x"00000010",
  1621 => x"00000000",
  1622 => x"13260000",
  1623 => x"00000000",
  1624 => x"00000000",
  1625 => x"00196900",
  1626 => x"4f4f4200",
  1627 => x"20202054",
  1628 => x"4d4f5220",
  1629 => x"f0fe1e00",
  1630 => x"cd78c048",
  1631 => x"26097909",
  1632 => x"fe1e1e4f",
  1633 => x"487ebff0",
  1634 => x"1e4f2626",
  1635 => x"c148f0fe",
  1636 => x"1e4f2678",
  1637 => x"c048f0fe",
  1638 => x"1e4f2678",
  1639 => x"52c04a71",
  1640 => x"0e4f2652",
  1641 => x"5d5c5b5e",
  1642 => x"7186f40e",
  1643 => x"7e6d974d",
  1644 => x"974ca5c1",
  1645 => x"a6c8486c",
  1646 => x"c4486e58",
  1647 => x"c505a866",
  1648 => x"c048ff87",
  1649 => x"caff87e6",
  1650 => x"49a5c287",
  1651 => x"714b6c97",
  1652 => x"6b974ba3",
  1653 => x"7e6c974b",
  1654 => x"80c1486e",
  1655 => x"c758a6c8",
  1656 => x"58a6cc98",
  1657 => x"fe7c9770",
  1658 => x"487387e1",
  1659 => x"4d268ef4",
  1660 => x"4b264c26",
  1661 => x"5e0e4f26",
  1662 => x"f40e5c5b",
  1663 => x"d84c7186",
  1664 => x"ffc34a66",
  1665 => x"4ba4c29a",
  1666 => x"73496c97",
  1667 => x"517249a1",
  1668 => x"6e7e6c97",
  1669 => x"c880c148",
  1670 => x"98c758a6",
  1671 => x"7058a6cc",
  1672 => x"ff8ef454",
  1673 => x"1e1e87ca",
  1674 => x"e087e8fd",
  1675 => x"c0494abf",
  1676 => x"0299c0e0",
  1677 => x"1e7287cb",
  1678 => x"49eeebc2",
  1679 => x"c487f7fe",
  1680 => x"87fdfc86",
  1681 => x"c2fd7e70",
  1682 => x"4f262687",
  1683 => x"eeebc21e",
  1684 => x"87c7fd49",
  1685 => x"49e6e8c1",
  1686 => x"c387dafc",
  1687 => x"4f2687f7",
  1688 => x"5c5b5e0e",
  1689 => x"4d710e5d",
  1690 => x"49eeebc2",
  1691 => x"7087f4fc",
  1692 => x"abb7c04b",
  1693 => x"87c2c304",
  1694 => x"05abf0c3",
  1695 => x"edc187c9",
  1696 => x"78c148c4",
  1697 => x"c387e3c2",
  1698 => x"c905abe0",
  1699 => x"c8edc187",
  1700 => x"c278c148",
  1701 => x"edc187d4",
  1702 => x"c602bfc8",
  1703 => x"a3c0c287",
  1704 => x"7387c24c",
  1705 => x"c4edc14c",
  1706 => x"e0c002bf",
  1707 => x"c4497487",
  1708 => x"c19129b7",
  1709 => x"7481e4ee",
  1710 => x"c29acf4a",
  1711 => x"7248c192",
  1712 => x"ff4a7030",
  1713 => x"694872ba",
  1714 => x"db797098",
  1715 => x"c4497487",
  1716 => x"c19129b7",
  1717 => x"7481e4ee",
  1718 => x"c29acf4a",
  1719 => x"7248c392",
  1720 => x"484a7030",
  1721 => x"7970b069",
  1722 => x"c0059d75",
  1723 => x"d0ff87f0",
  1724 => x"78e1c848",
  1725 => x"c548d4ff",
  1726 => x"c8edc178",
  1727 => x"87c302bf",
  1728 => x"c178e0c3",
  1729 => x"02bfc4ed",
  1730 => x"d4ff87c6",
  1731 => x"78f0c348",
  1732 => x"7b0bd4ff",
  1733 => x"48d0ff0b",
  1734 => x"c078e1c8",
  1735 => x"edc178e0",
  1736 => x"78c048c8",
  1737 => x"48c4edc1",
  1738 => x"ebc278c0",
  1739 => x"f2f949ee",
  1740 => x"c04b7087",
  1741 => x"fc03abb7",
  1742 => x"48c087fe",
  1743 => x"4c264d26",
  1744 => x"4f264b26",
  1745 => x"00000000",
  1746 => x"00000000",
  1747 => x"494a711e",
  1748 => x"2687cdfc",
  1749 => x"4ac01e4f",
  1750 => x"91c44972",
  1751 => x"81e4eec1",
  1752 => x"82c179c0",
  1753 => x"04aab7d0",
  1754 => x"4f2687ee",
  1755 => x"5c5b5e0e",
  1756 => x"4d710e5d",
  1757 => x"7587dcf8",
  1758 => x"2ab7c44a",
  1759 => x"e4eec192",
  1760 => x"cf4c7582",
  1761 => x"6a94c29c",
  1762 => x"2b744b49",
  1763 => x"48c29bc3",
  1764 => x"4c703074",
  1765 => x"4874bcff",
  1766 => x"7a709871",
  1767 => x"7387ecf7",
  1768 => x"87d8fe48",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"00000000",
  1776 => x"00000000",
  1777 => x"00000000",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"00000000",
  1783 => x"00000000",
  1784 => x"00000000",
  1785 => x"48d0ff1e",
  1786 => x"7178e1c8",
  1787 => x"08d4ff48",
  1788 => x"1e4f2678",
  1789 => x"c848d0ff",
  1790 => x"487178e1",
  1791 => x"7808d4ff",
  1792 => x"ff4866c4",
  1793 => x"267808d4",
  1794 => x"4a711e4f",
  1795 => x"1e4966c4",
  1796 => x"deff4972",
  1797 => x"48d0ff87",
  1798 => x"2678e0c0",
  1799 => x"731e4f26",
  1800 => x"c84b711e",
  1801 => x"731e4966",
  1802 => x"a2e0c14a",
  1803 => x"87d9ff49",
  1804 => x"2687c426",
  1805 => x"264c264d",
  1806 => x"1e4f264b",
  1807 => x"c34ad4ff",
  1808 => x"d0ff7aff",
  1809 => x"78e1c048",
  1810 => x"ebc27ade",
  1811 => x"497abff8",
  1812 => x"7028c848",
  1813 => x"d048717a",
  1814 => x"717a7028",
  1815 => x"7028d848",
  1816 => x"48d0ff7a",
  1817 => x"2678e0c0",
  1818 => x"d0ff1e4f",
  1819 => x"78c9c848",
  1820 => x"d4ff4871",
  1821 => x"4f267808",
  1822 => x"494a711e",
  1823 => x"d0ff87eb",
  1824 => x"2678c848",
  1825 => x"1e731e4f",
  1826 => x"ecc24b71",
  1827 => x"c302bfc8",
  1828 => x"87ebc287",
  1829 => x"c848d0ff",
  1830 => x"487378c9",
  1831 => x"ffb0e0c0",
  1832 => x"c27808d4",
  1833 => x"c048fceb",
  1834 => x"0266c878",
  1835 => x"ffc387c5",
  1836 => x"c087c249",
  1837 => x"c4ecc249",
  1838 => x"0266cc59",
  1839 => x"d5c587c6",
  1840 => x"87c44ad5",
  1841 => x"4affffcf",
  1842 => x"5ac8ecc2",
  1843 => x"48c8ecc2",
  1844 => x"87c478c1",
  1845 => x"4c264d26",
  1846 => x"4f264b26",
  1847 => x"5c5b5e0e",
  1848 => x"4a710e5d",
  1849 => x"bfc4ecc2",
  1850 => x"029a724c",
  1851 => x"c84987cb",
  1852 => x"fbf1c191",
  1853 => x"c483714b",
  1854 => x"fbf5c187",
  1855 => x"134dc04b",
  1856 => x"c2997449",
  1857 => x"48bfc0ec",
  1858 => x"d4ffb871",
  1859 => x"b7c17808",
  1860 => x"b7c8852c",
  1861 => x"87e704ad",
  1862 => x"bffcebc2",
  1863 => x"c280c848",
  1864 => x"fe58c0ec",
  1865 => x"731e87ee",
  1866 => x"134b711e",
  1867 => x"cb029a4a",
  1868 => x"fe497287",
  1869 => x"4a1387e6",
  1870 => x"87f5059a",
  1871 => x"1e87d9fe",
  1872 => x"bffcebc2",
  1873 => x"fcebc249",
  1874 => x"78a1c148",
  1875 => x"a9b7c0c4",
  1876 => x"ff87db03",
  1877 => x"ecc248d4",
  1878 => x"c278bfc0",
  1879 => x"49bffceb",
  1880 => x"48fcebc2",
  1881 => x"c478a1c1",
  1882 => x"04a9b7c0",
  1883 => x"d0ff87e5",
  1884 => x"c278c848",
  1885 => x"c048c8ec",
  1886 => x"004f2678",
  1887 => x"00000000",
  1888 => x"00000000",
  1889 => x"5f5f0000",
  1890 => x"00000000",
  1891 => x"03000303",
  1892 => x"14000003",
  1893 => x"7f147f7f",
  1894 => x"0000147f",
  1895 => x"6b6b2e24",
  1896 => x"4c00123a",
  1897 => x"6c18366a",
  1898 => x"30003256",
  1899 => x"77594f7e",
  1900 => x"0040683a",
  1901 => x"03070400",
  1902 => x"00000000",
  1903 => x"633e1c00",
  1904 => x"00000041",
  1905 => x"3e634100",
  1906 => x"0800001c",
  1907 => x"1c1c3e2a",
  1908 => x"00082a3e",
  1909 => x"3e3e0808",
  1910 => x"00000808",
  1911 => x"60e08000",
  1912 => x"00000000",
  1913 => x"08080808",
  1914 => x"00000808",
  1915 => x"60600000",
  1916 => x"40000000",
  1917 => x"0c183060",
  1918 => x"00010306",
  1919 => x"4d597f3e",
  1920 => x"00003e7f",
  1921 => x"7f7f0604",
  1922 => x"00000000",
  1923 => x"59716342",
  1924 => x"0000464f",
  1925 => x"49496322",
  1926 => x"1800367f",
  1927 => x"7f13161c",
  1928 => x"0000107f",
  1929 => x"45456727",
  1930 => x"0000397d",
  1931 => x"494b7e3c",
  1932 => x"00003079",
  1933 => x"79710101",
  1934 => x"0000070f",
  1935 => x"49497f36",
  1936 => x"0000367f",
  1937 => x"69494f06",
  1938 => x"00001e3f",
  1939 => x"66660000",
  1940 => x"00000000",
  1941 => x"66e68000",
  1942 => x"00000000",
  1943 => x"14140808",
  1944 => x"00002222",
  1945 => x"14141414",
  1946 => x"00001414",
  1947 => x"14142222",
  1948 => x"00000808",
  1949 => x"59510302",
  1950 => x"3e00060f",
  1951 => x"555d417f",
  1952 => x"00001e1f",
  1953 => x"09097f7e",
  1954 => x"00007e7f",
  1955 => x"49497f7f",
  1956 => x"0000367f",
  1957 => x"41633e1c",
  1958 => x"00004141",
  1959 => x"63417f7f",
  1960 => x"00001c3e",
  1961 => x"49497f7f",
  1962 => x"00004141",
  1963 => x"09097f7f",
  1964 => x"00000101",
  1965 => x"49417f3e",
  1966 => x"00007a7b",
  1967 => x"08087f7f",
  1968 => x"00007f7f",
  1969 => x"7f7f4100",
  1970 => x"00000041",
  1971 => x"40406020",
  1972 => x"7f003f7f",
  1973 => x"361c087f",
  1974 => x"00004163",
  1975 => x"40407f7f",
  1976 => x"7f004040",
  1977 => x"060c067f",
  1978 => x"7f007f7f",
  1979 => x"180c067f",
  1980 => x"00007f7f",
  1981 => x"41417f3e",
  1982 => x"00003e7f",
  1983 => x"09097f7f",
  1984 => x"3e00060f",
  1985 => x"7f61417f",
  1986 => x"0000407e",
  1987 => x"19097f7f",
  1988 => x"0000667f",
  1989 => x"594d6f26",
  1990 => x"0000327b",
  1991 => x"7f7f0101",
  1992 => x"00000101",
  1993 => x"40407f3f",
  1994 => x"00003f7f",
  1995 => x"70703f0f",
  1996 => x"7f000f3f",
  1997 => x"3018307f",
  1998 => x"41007f7f",
  1999 => x"1c1c3663",
  2000 => x"01416336",
  2001 => x"7c7c0603",
  2002 => x"61010306",
  2003 => x"474d5971",
  2004 => x"00004143",
  2005 => x"417f7f00",
  2006 => x"01000041",
  2007 => x"180c0603",
  2008 => x"00406030",
  2009 => x"7f414100",
  2010 => x"0800007f",
  2011 => x"0603060c",
  2012 => x"8000080c",
  2013 => x"80808080",
  2014 => x"00008080",
  2015 => x"07030000",
  2016 => x"00000004",
  2017 => x"54547420",
  2018 => x"0000787c",
  2019 => x"44447f7f",
  2020 => x"0000387c",
  2021 => x"44447c38",
  2022 => x"00000044",
  2023 => x"44447c38",
  2024 => x"00007f7f",
  2025 => x"54547c38",
  2026 => x"0000185c",
  2027 => x"057f7e04",
  2028 => x"00000005",
  2029 => x"a4a4bc18",
  2030 => x"00007cfc",
  2031 => x"04047f7f",
  2032 => x"0000787c",
  2033 => x"7d3d0000",
  2034 => x"00000040",
  2035 => x"fd808080",
  2036 => x"0000007d",
  2037 => x"38107f7f",
  2038 => x"0000446c",
  2039 => x"7f3f0000",
  2040 => x"7c000040",
  2041 => x"0c180c7c",
  2042 => x"0000787c",
  2043 => x"04047c7c",
  2044 => x"0000787c",
  2045 => x"44447c38",
  2046 => x"0000387c",
  2047 => x"2424fcfc",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
