library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0000183c",
     1 => x"24243c18",
     2 => x"0000fcfc",
     3 => x"04047c7c",
     4 => x"0000080c",
     5 => x"54545c48",
     6 => x"00002074",
     7 => x"447f3f04",
     8 => x"00000044",
     9 => x"40407c3c",
    10 => x"00007c7c",
    11 => x"60603c1c",
    12 => x"3c001c3c",
    13 => x"6030607c",
    14 => x"44003c7c",
    15 => x"3810386c",
    16 => x"0000446c",
    17 => x"60e0bc1c",
    18 => x"00001c3c",
    19 => x"5c746444",
    20 => x"0000444c",
    21 => x"773e0808",
    22 => x"00004141",
    23 => x"7f7f0000",
    24 => x"00000000",
    25 => x"3e774141",
    26 => x"02000808",
    27 => x"02030101",
    28 => x"7f000102",
    29 => x"7f7f7f7f",
    30 => x"08007f7f",
    31 => x"3e1c1c08",
    32 => x"7f7f7f3e",
    33 => x"1c3e3e7f",
    34 => x"0008081c",
    35 => x"7c7c1810",
    36 => x"00001018",
    37 => x"7c7c3010",
    38 => x"10001030",
    39 => x"78606030",
    40 => x"4200061e",
    41 => x"3c183c66",
    42 => x"78004266",
    43 => x"c6c26a38",
    44 => x"6000386c",
    45 => x"00600000",
    46 => x"0e006000",
    47 => x"5d5c5b5e",
    48 => x"4c711e0e",
    49 => x"bfd9ecc2",
    50 => x"c04bc04d",
    51 => x"02ab741e",
    52 => x"a6c487c7",
    53 => x"c578c048",
    54 => x"48a6c487",
    55 => x"66c478c1",
    56 => x"ee49731e",
    57 => x"86c887df",
    58 => x"ef49e0c0",
    59 => x"a5c487ee",
    60 => x"f0496a4a",
    61 => x"c6f187f0",
    62 => x"c185cb87",
    63 => x"abb7c883",
    64 => x"87c7ff04",
    65 => x"264d2626",
    66 => x"264b264c",
    67 => x"4a711e4f",
    68 => x"5addecc2",
    69 => x"48ddecc2",
    70 => x"fe4978c7",
    71 => x"4f2687dd",
    72 => x"711e731e",
    73 => x"aab7c04a",
    74 => x"c287d303",
    75 => x"05bfdcd2",
    76 => x"4bc187c4",
    77 => x"4bc087c2",
    78 => x"5be0d2c2",
    79 => x"d2c287c4",
    80 => x"d2c25ae0",
    81 => x"c14abfdc",
    82 => x"a2c0c19a",
    83 => x"87e8ec49",
    84 => x"d2c248fc",
    85 => x"fe78bfdc",
    86 => x"711e87ef",
    87 => x"1e66c44a",
    88 => x"f9ea4972",
    89 => x"4f262687",
    90 => x"48d4ff1e",
    91 => x"ff78ffc3",
    92 => x"e1c048d0",
    93 => x"48d4ff78",
    94 => x"487178c1",
    95 => x"d4ff30c4",
    96 => x"d0ff7808",
    97 => x"78e0c048",
    98 => x"c21e4f26",
    99 => x"49bfdcd2",
   100 => x"c287f9e6",
   101 => x"e848d1ec",
   102 => x"ecc278bf",
   103 => x"bfec48cd",
   104 => x"d1ecc278",
   105 => x"c3494abf",
   106 => x"b7c899ff",
   107 => x"7148722a",
   108 => x"d9ecc2b0",
   109 => x"0e4f2658",
   110 => x"5d5c5b5e",
   111 => x"ff4b710e",
   112 => x"ecc287c8",
   113 => x"50c048cc",
   114 => x"dfe64973",
   115 => x"4c497087",
   116 => x"eecb9cc2",
   117 => x"87cccb49",
   118 => x"ecc24d70",
   119 => x"05bf97cc",
   120 => x"d087e2c1",
   121 => x"ecc24966",
   122 => x"0599bfd5",
   123 => x"66d487d6",
   124 => x"cdecc249",
   125 => x"cb0599bf",
   126 => x"e5497387",
   127 => x"987087ee",
   128 => x"87c1c102",
   129 => x"c1fe4cc1",
   130 => x"ca497587",
   131 => x"987087e2",
   132 => x"c287c602",
   133 => x"c148ccec",
   134 => x"ccecc250",
   135 => x"c005bf97",
   136 => x"ecc287e3",
   137 => x"d049bfd5",
   138 => x"ff059966",
   139 => x"ecc287d6",
   140 => x"d449bfcd",
   141 => x"ff059966",
   142 => x"497387ca",
   143 => x"7087ede4",
   144 => x"fffe0598",
   145 => x"fa487487",
   146 => x"5e0e87fb",
   147 => x"0e5d5c5b",
   148 => x"4dc086f8",
   149 => x"7ebfec4c",
   150 => x"c248a6c4",
   151 => x"78bfd9ec",
   152 => x"1ec01ec1",
   153 => x"cefd49c7",
   154 => x"7086c887",
   155 => x"87cd0298",
   156 => x"ebfa49ff",
   157 => x"49dac187",
   158 => x"c187f1e3",
   159 => x"ccecc24d",
   160 => x"cf02bf97",
   161 => x"d4d2c287",
   162 => x"b9c149bf",
   163 => x"59d8d2c2",
   164 => x"87d4fb71",
   165 => x"bfd1ecc2",
   166 => x"dcd2c24b",
   167 => x"e9c005bf",
   168 => x"49fdc387",
   169 => x"c387c5e3",
   170 => x"ffe249fa",
   171 => x"c3497387",
   172 => x"1e7199ff",
   173 => x"e1fa49c0",
   174 => x"c8497387",
   175 => x"1e7129b7",
   176 => x"d5fa49c1",
   177 => x"c586c887",
   178 => x"ecc287f4",
   179 => x"9b4bbfd5",
   180 => x"c287dd02",
   181 => x"49bfd8d2",
   182 => x"7087d5c7",
   183 => x"87c40598",
   184 => x"87d24bc0",
   185 => x"c649e0c2",
   186 => x"d2c287fa",
   187 => x"87c658dc",
   188 => x"48d8d2c2",
   189 => x"497378c0",
   190 => x"cd0599c2",
   191 => x"49ebc387",
   192 => x"7087e9e1",
   193 => x"0299c249",
   194 => x"4cfb87c2",
   195 => x"99c14973",
   196 => x"c387cd05",
   197 => x"d3e149f4",
   198 => x"c2497087",
   199 => x"87c20299",
   200 => x"49734cfa",
   201 => x"cd0599c8",
   202 => x"49f5c387",
   203 => x"7087fde0",
   204 => x"0299c249",
   205 => x"ecc287d5",
   206 => x"ca02bfdd",
   207 => x"88c14887",
   208 => x"58e1ecc2",
   209 => x"ff87c2c0",
   210 => x"734dc14c",
   211 => x"0599c449",
   212 => x"f2c387cd",
   213 => x"87d4e049",
   214 => x"99c24970",
   215 => x"c287dc02",
   216 => x"7ebfddec",
   217 => x"a8b7c748",
   218 => x"87cbc003",
   219 => x"80c1486e",
   220 => x"58e1ecc2",
   221 => x"fe87c2c0",
   222 => x"c34dc14c",
   223 => x"dfff49fd",
   224 => x"497087ea",
   225 => x"d50299c2",
   226 => x"ddecc287",
   227 => x"c9c002bf",
   228 => x"ddecc287",
   229 => x"c078c048",
   230 => x"4cfd87c2",
   231 => x"fac34dc1",
   232 => x"c7dfff49",
   233 => x"c2497087",
   234 => x"d9c00299",
   235 => x"ddecc287",
   236 => x"b7c748bf",
   237 => x"c9c003a8",
   238 => x"ddecc287",
   239 => x"c078c748",
   240 => x"4cfc87c2",
   241 => x"b7c04dc1",
   242 => x"d3c003ac",
   243 => x"4866c487",
   244 => x"7080d8c1",
   245 => x"02bf6e7e",
   246 => x"4b87c5c0",
   247 => x"0f734974",
   248 => x"f0c31ec0",
   249 => x"49dac11e",
   250 => x"c887ccf7",
   251 => x"02987086",
   252 => x"c287d8c0",
   253 => x"7ebfddec",
   254 => x"91cb496e",
   255 => x"714a66c4",
   256 => x"c0026a82",
   257 => x"6e4b87c5",
   258 => x"750f7349",
   259 => x"c8c0029d",
   260 => x"ddecc287",
   261 => x"e2f249bf",
   262 => x"e0d2c287",
   263 => x"ddc002bf",
   264 => x"cbc24987",
   265 => x"02987087",
   266 => x"c287d3c0",
   267 => x"49bfddec",
   268 => x"c087c8f2",
   269 => x"87e8f349",
   270 => x"48e0d2c2",
   271 => x"8ef878c0",
   272 => x"0e87c2f3",
   273 => x"5d5c5b5e",
   274 => x"4c711e0e",
   275 => x"bfd9ecc2",
   276 => x"a1cdc149",
   277 => x"81d1c14d",
   278 => x"9c747e69",
   279 => x"c487cf02",
   280 => x"7b744ba5",
   281 => x"bfd9ecc2",
   282 => x"87e1f249",
   283 => x"9c747b6e",
   284 => x"c087c405",
   285 => x"c187c24b",
   286 => x"f249734b",
   287 => x"66d487e2",
   288 => x"4987c702",
   289 => x"4a7087de",
   290 => x"4ac087c2",
   291 => x"5ae4d2c2",
   292 => x"87f1f126",
   293 => x"00000000",
   294 => x"00000000",
   295 => x"00000000",
   296 => x"00000000",
   297 => x"ff4a711e",
   298 => x"7249bfc8",
   299 => x"4f2648a1",
   300 => x"bfc8ff1e",
   301 => x"c0c0fe89",
   302 => x"a9c0c0c0",
   303 => x"c087c401",
   304 => x"c187c24a",
   305 => x"2648724a",
   306 => x"5b5e0e4f",
   307 => x"710e5d5c",
   308 => x"4cd4ff4b",
   309 => x"c04866d0",
   310 => x"ff49d678",
   311 => x"c387c5dc",
   312 => x"496c7cff",
   313 => x"7199ffc3",
   314 => x"f0c3494d",
   315 => x"a9e0c199",
   316 => x"c387cb05",
   317 => x"486c7cff",
   318 => x"66d098c3",
   319 => x"ffc37808",
   320 => x"494a6c7c",
   321 => x"ffc331c8",
   322 => x"714a6c7c",
   323 => x"c84972b2",
   324 => x"7cffc331",
   325 => x"b2714a6c",
   326 => x"31c84972",
   327 => x"6c7cffc3",
   328 => x"ffb2714a",
   329 => x"e0c048d0",
   330 => x"029b7378",
   331 => x"7b7287c2",
   332 => x"4d264875",
   333 => x"4b264c26",
   334 => x"261e4f26",
   335 => x"5b5e0e4f",
   336 => x"86f80e5c",
   337 => x"a6c81e76",
   338 => x"87fdfd49",
   339 => x"4b7086c4",
   340 => x"a8c8486e",
   341 => x"87f0c203",
   342 => x"f0c34a73",
   343 => x"aad0c19a",
   344 => x"c187c702",
   345 => x"c205aae0",
   346 => x"497387de",
   347 => x"c30299c8",
   348 => x"87c6ff87",
   349 => x"9cc34c73",
   350 => x"c105acc2",
   351 => x"66c487c2",
   352 => x"7131c949",
   353 => x"4a66c41e",
   354 => x"ecc292d4",
   355 => x"817249e1",
   356 => x"87f3d0fe",
   357 => x"d9ff49d8",
   358 => x"c0c887ca",
   359 => x"fedac21e",
   360 => x"f9ecfd49",
   361 => x"48d0ff87",
   362 => x"c278e0c0",
   363 => x"cc1efeda",
   364 => x"92d44a66",
   365 => x"49e1ecc2",
   366 => x"cefe8172",
   367 => x"86cc87fb",
   368 => x"c105acc1",
   369 => x"66c487c2",
   370 => x"7131c949",
   371 => x"4a66c41e",
   372 => x"ecc292d4",
   373 => x"817249e1",
   374 => x"87ebcffe",
   375 => x"1efedac2",
   376 => x"d44a66c8",
   377 => x"e1ecc292",
   378 => x"fe817249",
   379 => x"d787fccc",
   380 => x"efd7ff49",
   381 => x"1ec0c887",
   382 => x"49fedac2",
   383 => x"87f7eafd",
   384 => x"d0ff86cc",
   385 => x"78e0c048",
   386 => x"e7fc8ef8",
   387 => x"5b5e0e87",
   388 => x"1e0e5d5c",
   389 => x"d4ff4d71",
   390 => x"7e66d44c",
   391 => x"a8b7c348",
   392 => x"c087c506",
   393 => x"87e9c148",
   394 => x"ddfe4975",
   395 => x"1e7587e0",
   396 => x"d44b66c4",
   397 => x"e1ecc293",
   398 => x"fe497383",
   399 => x"c887fac6",
   400 => x"ff4b6b83",
   401 => x"e1c848d0",
   402 => x"737cdd78",
   403 => x"98ffc348",
   404 => x"49737c70",
   405 => x"7129b7c8",
   406 => x"98ffc348",
   407 => x"49737c70",
   408 => x"7129b7d0",
   409 => x"98ffc348",
   410 => x"48737c70",
   411 => x"7028b7d8",
   412 => x"7c7cc07c",
   413 => x"7c7c7c7c",
   414 => x"7c7c7c7c",
   415 => x"d0ff7c7c",
   416 => x"78e0c048",
   417 => x"dc1e66c4",
   418 => x"fcd5ff49",
   419 => x"7386c887",
   420 => x"ddfa2648",
   421 => x"ddfa2687",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
