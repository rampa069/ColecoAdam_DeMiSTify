
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"c4",x"ef",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"c4",x"ef",x"c2"),
    14 => (x"48",x"d8",x"da",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"cd",x"e2"),
    19 => (x"72",x"1e",x"87",x"fd"),
    20 => (x"12",x"1e",x"73",x"1e"),
    21 => (x"ca",x"02",x"11",x"48"),
    22 => (x"df",x"c3",x"4b",x"87"),
    23 => (x"88",x"73",x"9b",x"98"),
    24 => (x"26",x"87",x"f0",x"02"),
    25 => (x"26",x"4a",x"26",x"4b"),
    26 => (x"1e",x"73",x"1e",x"4f"),
    27 => (x"8b",x"c1",x"1e",x"72"),
    28 => (x"12",x"87",x"ca",x"04"),
    29 => (x"c4",x"02",x"11",x"48"),
    30 => (x"f1",x"02",x"88",x"87"),
    31 => (x"26",x"4a",x"26",x"87"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"1e",x"73",x"1e",x"74"),
    34 => (x"8b",x"c1",x"1e",x"72"),
    35 => (x"12",x"87",x"d0",x"04"),
    36 => (x"ca",x"02",x"11",x"48"),
    37 => (x"df",x"c3",x"4c",x"87"),
    38 => (x"88",x"74",x"9c",x"98"),
    39 => (x"26",x"87",x"eb",x"02"),
    40 => (x"26",x"4b",x"26",x"4a"),
    41 => (x"1e",x"4f",x"26",x"4c"),
    42 => (x"73",x"81",x"48",x"73"),
    43 => (x"87",x"c5",x"02",x"a9"),
    44 => (x"f6",x"05",x"53",x"12"),
    45 => (x"1e",x"4f",x"26",x"87"),
    46 => (x"66",x"c4",x"4a",x"71"),
    47 => (x"88",x"c1",x"48",x"49"),
    48 => (x"71",x"58",x"a6",x"c8"),
    49 => (x"87",x"d4",x"02",x"99"),
    50 => (x"d4",x"ff",x"48",x"12"),
    51 => (x"66",x"c4",x"78",x"08"),
    52 => (x"88",x"c1",x"48",x"49"),
    53 => (x"71",x"58",x"a6",x"c8"),
    54 => (x"87",x"ec",x"05",x"99"),
    55 => (x"71",x"1e",x"4f",x"26"),
    56 => (x"49",x"66",x"c4",x"4a"),
    57 => (x"c8",x"88",x"c1",x"48"),
    58 => (x"99",x"71",x"58",x"a6"),
    59 => (x"ff",x"87",x"d6",x"02"),
    60 => (x"ff",x"c3",x"48",x"d4"),
    61 => (x"c4",x"52",x"68",x"78"),
    62 => (x"c1",x"48",x"49",x"66"),
    63 => (x"58",x"a6",x"c8",x"88"),
    64 => (x"ea",x"05",x"99",x"71"),
    65 => (x"1e",x"4f",x"26",x"87"),
    66 => (x"d4",x"ff",x"1e",x"73"),
    67 => (x"7b",x"ff",x"c3",x"4b"),
    68 => (x"ff",x"c3",x"4a",x"6b"),
    69 => (x"c8",x"49",x"6b",x"7b"),
    70 => (x"c3",x"b1",x"72",x"32"),
    71 => (x"4a",x"6b",x"7b",x"ff"),
    72 => (x"b2",x"71",x"31",x"c8"),
    73 => (x"6b",x"7b",x"ff",x"c3"),
    74 => (x"72",x"32",x"c8",x"49"),
    75 => (x"c4",x"48",x"71",x"b1"),
    76 => (x"26",x"4d",x"26",x"87"),
    77 => (x"26",x"4b",x"26",x"4c"),
    78 => (x"5b",x"5e",x"0e",x"4f"),
    79 => (x"71",x"0e",x"5d",x"5c"),
    80 => (x"4c",x"d4",x"ff",x"4a"),
    81 => (x"ff",x"c3",x"48",x"72"),
    82 => (x"c2",x"7c",x"70",x"98"),
    83 => (x"05",x"bf",x"d8",x"da"),
    84 => (x"66",x"d0",x"87",x"c8"),
    85 => (x"d4",x"30",x"c9",x"48"),
    86 => (x"66",x"d0",x"58",x"a6"),
    87 => (x"71",x"29",x"d8",x"49"),
    88 => (x"98",x"ff",x"c3",x"48"),
    89 => (x"66",x"d0",x"7c",x"70"),
    90 => (x"71",x"29",x"d0",x"49"),
    91 => (x"98",x"ff",x"c3",x"48"),
    92 => (x"66",x"d0",x"7c",x"70"),
    93 => (x"71",x"29",x"c8",x"49"),
    94 => (x"98",x"ff",x"c3",x"48"),
    95 => (x"66",x"d0",x"7c",x"70"),
    96 => (x"98",x"ff",x"c3",x"48"),
    97 => (x"49",x"72",x"7c",x"70"),
    98 => (x"48",x"71",x"29",x"d0"),
    99 => (x"70",x"98",x"ff",x"c3"),
   100 => (x"c9",x"4b",x"6c",x"7c"),
   101 => (x"c3",x"4d",x"ff",x"f0"),
   102 => (x"d0",x"05",x"ab",x"ff"),
   103 => (x"7c",x"ff",x"c3",x"87"),
   104 => (x"8d",x"c1",x"4b",x"6c"),
   105 => (x"c3",x"87",x"c6",x"02"),
   106 => (x"f0",x"02",x"ab",x"ff"),
   107 => (x"fd",x"48",x"73",x"87"),
   108 => (x"c0",x"1e",x"87",x"ff"),
   109 => (x"48",x"d4",x"ff",x"49"),
   110 => (x"c1",x"78",x"ff",x"c3"),
   111 => (x"b7",x"c8",x"c3",x"81"),
   112 => (x"87",x"f1",x"04",x"a9"),
   113 => (x"73",x"1e",x"4f",x"26"),
   114 => (x"c4",x"87",x"e7",x"1e"),
   115 => (x"c0",x"4b",x"df",x"f8"),
   116 => (x"f0",x"ff",x"c0",x"1e"),
   117 => (x"fd",x"49",x"f7",x"c1"),
   118 => (x"86",x"c4",x"87",x"df"),
   119 => (x"c0",x"05",x"a8",x"c1"),
   120 => (x"d4",x"ff",x"87",x"ea"),
   121 => (x"78",x"ff",x"c3",x"48"),
   122 => (x"c0",x"c0",x"c0",x"c1"),
   123 => (x"c0",x"1e",x"c0",x"c0"),
   124 => (x"e9",x"c1",x"f0",x"e1"),
   125 => (x"87",x"c1",x"fd",x"49"),
   126 => (x"98",x"70",x"86",x"c4"),
   127 => (x"ff",x"87",x"ca",x"05"),
   128 => (x"ff",x"c3",x"48",x"d4"),
   129 => (x"cb",x"48",x"c1",x"78"),
   130 => (x"87",x"e6",x"fe",x"87"),
   131 => (x"fe",x"05",x"8b",x"c1"),
   132 => (x"48",x"c0",x"87",x"fd"),
   133 => (x"1e",x"87",x"de",x"fc"),
   134 => (x"d4",x"ff",x"1e",x"73"),
   135 => (x"78",x"ff",x"c3",x"48"),
   136 => (x"1e",x"c0",x"4b",x"d3"),
   137 => (x"c1",x"f0",x"ff",x"c0"),
   138 => (x"cc",x"fc",x"49",x"c1"),
   139 => (x"70",x"86",x"c4",x"87"),
   140 => (x"87",x"ca",x"05",x"98"),
   141 => (x"c3",x"48",x"d4",x"ff"),
   142 => (x"48",x"c1",x"78",x"ff"),
   143 => (x"f1",x"fd",x"87",x"cb"),
   144 => (x"05",x"8b",x"c1",x"87"),
   145 => (x"c0",x"87",x"db",x"ff"),
   146 => (x"87",x"e9",x"fb",x"48"),
   147 => (x"5c",x"5b",x"5e",x"0e"),
   148 => (x"4c",x"d4",x"ff",x"0e"),
   149 => (x"c6",x"87",x"db",x"fd"),
   150 => (x"e1",x"c0",x"1e",x"ea"),
   151 => (x"49",x"c8",x"c1",x"f0"),
   152 => (x"c4",x"87",x"d6",x"fb"),
   153 => (x"02",x"a8",x"c1",x"86"),
   154 => (x"ea",x"fe",x"87",x"c8"),
   155 => (x"c1",x"48",x"c0",x"87"),
   156 => (x"d2",x"fa",x"87",x"e2"),
   157 => (x"cf",x"49",x"70",x"87"),
   158 => (x"c6",x"99",x"ff",x"ff"),
   159 => (x"c8",x"02",x"a9",x"ea"),
   160 => (x"87",x"d3",x"fe",x"87"),
   161 => (x"cb",x"c1",x"48",x"c0"),
   162 => (x"7c",x"ff",x"c3",x"87"),
   163 => (x"fc",x"4b",x"f1",x"c0"),
   164 => (x"98",x"70",x"87",x"f4"),
   165 => (x"87",x"eb",x"c0",x"02"),
   166 => (x"ff",x"c0",x"1e",x"c0"),
   167 => (x"49",x"fa",x"c1",x"f0"),
   168 => (x"c4",x"87",x"d6",x"fa"),
   169 => (x"05",x"98",x"70",x"86"),
   170 => (x"ff",x"c3",x"87",x"d9"),
   171 => (x"c3",x"49",x"6c",x"7c"),
   172 => (x"7c",x"7c",x"7c",x"ff"),
   173 => (x"99",x"c0",x"c1",x"7c"),
   174 => (x"c1",x"87",x"c4",x"02"),
   175 => (x"c0",x"87",x"d5",x"48"),
   176 => (x"c2",x"87",x"d1",x"48"),
   177 => (x"87",x"c4",x"05",x"ab"),
   178 => (x"87",x"c8",x"48",x"c0"),
   179 => (x"fe",x"05",x"8b",x"c1"),
   180 => (x"48",x"c0",x"87",x"fd"),
   181 => (x"1e",x"87",x"dc",x"f9"),
   182 => (x"da",x"c2",x"1e",x"73"),
   183 => (x"78",x"c1",x"48",x"d8"),
   184 => (x"d0",x"ff",x"4b",x"c7"),
   185 => (x"fb",x"78",x"c2",x"48"),
   186 => (x"d0",x"ff",x"87",x"c8"),
   187 => (x"c0",x"78",x"c3",x"48"),
   188 => (x"d0",x"e5",x"c0",x"1e"),
   189 => (x"f8",x"49",x"c0",x"c1"),
   190 => (x"86",x"c4",x"87",x"ff"),
   191 => (x"c1",x"05",x"a8",x"c1"),
   192 => (x"ab",x"c2",x"4b",x"87"),
   193 => (x"c0",x"87",x"c5",x"05"),
   194 => (x"87",x"f9",x"c0",x"48"),
   195 => (x"ff",x"05",x"8b",x"c1"),
   196 => (x"f7",x"fc",x"87",x"d0"),
   197 => (x"dc",x"da",x"c2",x"87"),
   198 => (x"05",x"98",x"70",x"58"),
   199 => (x"1e",x"c1",x"87",x"cd"),
   200 => (x"c1",x"f0",x"ff",x"c0"),
   201 => (x"d0",x"f8",x"49",x"d0"),
   202 => (x"ff",x"86",x"c4",x"87"),
   203 => (x"ff",x"c3",x"48",x"d4"),
   204 => (x"87",x"dd",x"c4",x"78"),
   205 => (x"58",x"e0",x"da",x"c2"),
   206 => (x"c2",x"48",x"d0",x"ff"),
   207 => (x"48",x"d4",x"ff",x"78"),
   208 => (x"c1",x"78",x"ff",x"c3"),
   209 => (x"87",x"ed",x"f7",x"48"),
   210 => (x"5c",x"5b",x"5e",x"0e"),
   211 => (x"4a",x"71",x"0e",x"5d"),
   212 => (x"ff",x"4d",x"ff",x"c3"),
   213 => (x"7c",x"75",x"4c",x"d4"),
   214 => (x"c4",x"48",x"d0",x"ff"),
   215 => (x"7c",x"75",x"78",x"c3"),
   216 => (x"ff",x"c0",x"1e",x"72"),
   217 => (x"49",x"d8",x"c1",x"f0"),
   218 => (x"c4",x"87",x"ce",x"f7"),
   219 => (x"02",x"98",x"70",x"86"),
   220 => (x"48",x"c1",x"87",x"c5"),
   221 => (x"75",x"87",x"ee",x"c0"),
   222 => (x"7c",x"fe",x"c3",x"7c"),
   223 => (x"d4",x"1e",x"c0",x"c8"),
   224 => (x"f2",x"f4",x"49",x"66"),
   225 => (x"75",x"86",x"c4",x"87"),
   226 => (x"75",x"7c",x"75",x"7c"),
   227 => (x"e0",x"da",x"d8",x"7c"),
   228 => (x"6c",x"7c",x"75",x"4b"),
   229 => (x"c1",x"87",x"c5",x"05"),
   230 => (x"87",x"f5",x"05",x"8b"),
   231 => (x"d0",x"ff",x"7c",x"75"),
   232 => (x"c0",x"78",x"c2",x"48"),
   233 => (x"87",x"c9",x"f6",x"48"),
   234 => (x"5c",x"5b",x"5e",x"0e"),
   235 => (x"4b",x"71",x"0e",x"5d"),
   236 => (x"ee",x"c5",x"4c",x"c0"),
   237 => (x"ff",x"4a",x"df",x"cd"),
   238 => (x"ff",x"c3",x"48",x"d4"),
   239 => (x"c3",x"48",x"68",x"78"),
   240 => (x"c0",x"05",x"a8",x"fe"),
   241 => (x"d4",x"ff",x"87",x"fe"),
   242 => (x"02",x"9b",x"73",x"4d"),
   243 => (x"66",x"d0",x"87",x"cc"),
   244 => (x"f4",x"49",x"73",x"1e"),
   245 => (x"86",x"c4",x"87",x"c8"),
   246 => (x"d0",x"ff",x"87",x"d6"),
   247 => (x"78",x"d1",x"c4",x"48"),
   248 => (x"d0",x"7d",x"ff",x"c3"),
   249 => (x"88",x"c1",x"48",x"66"),
   250 => (x"70",x"58",x"a6",x"d4"),
   251 => (x"87",x"f0",x"05",x"98"),
   252 => (x"c3",x"48",x"d4",x"ff"),
   253 => (x"73",x"78",x"78",x"ff"),
   254 => (x"87",x"c5",x"05",x"9b"),
   255 => (x"d0",x"48",x"d0",x"ff"),
   256 => (x"4c",x"4a",x"c1",x"78"),
   257 => (x"fe",x"05",x"8a",x"c1"),
   258 => (x"48",x"74",x"87",x"ed"),
   259 => (x"1e",x"87",x"e2",x"f4"),
   260 => (x"4a",x"71",x"1e",x"73"),
   261 => (x"d4",x"ff",x"4b",x"c0"),
   262 => (x"78",x"ff",x"c3",x"48"),
   263 => (x"c4",x"48",x"d0",x"ff"),
   264 => (x"d4",x"ff",x"78",x"c3"),
   265 => (x"78",x"ff",x"c3",x"48"),
   266 => (x"ff",x"c0",x"1e",x"72"),
   267 => (x"49",x"d1",x"c1",x"f0"),
   268 => (x"c4",x"87",x"c6",x"f4"),
   269 => (x"05",x"98",x"70",x"86"),
   270 => (x"c0",x"c8",x"87",x"d2"),
   271 => (x"49",x"66",x"cc",x"1e"),
   272 => (x"c4",x"87",x"e5",x"fd"),
   273 => (x"ff",x"4b",x"70",x"86"),
   274 => (x"78",x"c2",x"48",x"d0"),
   275 => (x"e4",x"f3",x"48",x"73"),
   276 => (x"5b",x"5e",x"0e",x"87"),
   277 => (x"c0",x"0e",x"5d",x"5c"),
   278 => (x"f0",x"ff",x"c0",x"1e"),
   279 => (x"f3",x"49",x"c9",x"c1"),
   280 => (x"1e",x"d2",x"87",x"d7"),
   281 => (x"49",x"e0",x"da",x"c2"),
   282 => (x"c8",x"87",x"fd",x"fc"),
   283 => (x"c1",x"4c",x"c0",x"86"),
   284 => (x"ac",x"b7",x"d2",x"84"),
   285 => (x"c2",x"87",x"f8",x"04"),
   286 => (x"bf",x"97",x"e0",x"da"),
   287 => (x"99",x"c0",x"c3",x"49"),
   288 => (x"05",x"a9",x"c0",x"c1"),
   289 => (x"c2",x"87",x"e7",x"c0"),
   290 => (x"bf",x"97",x"e7",x"da"),
   291 => (x"c2",x"31",x"d0",x"49"),
   292 => (x"bf",x"97",x"e8",x"da"),
   293 => (x"72",x"32",x"c8",x"4a"),
   294 => (x"e9",x"da",x"c2",x"b1"),
   295 => (x"b1",x"4a",x"bf",x"97"),
   296 => (x"ff",x"cf",x"4c",x"71"),
   297 => (x"c1",x"9c",x"ff",x"ff"),
   298 => (x"c1",x"34",x"ca",x"84"),
   299 => (x"da",x"c2",x"87",x"e7"),
   300 => (x"49",x"bf",x"97",x"e9"),
   301 => (x"99",x"c6",x"31",x"c1"),
   302 => (x"97",x"ea",x"da",x"c2"),
   303 => (x"b7",x"c7",x"4a",x"bf"),
   304 => (x"c2",x"b1",x"72",x"2a"),
   305 => (x"bf",x"97",x"e5",x"da"),
   306 => (x"9d",x"cf",x"4d",x"4a"),
   307 => (x"97",x"e6",x"da",x"c2"),
   308 => (x"9a",x"c3",x"4a",x"bf"),
   309 => (x"da",x"c2",x"32",x"ca"),
   310 => (x"4b",x"bf",x"97",x"e7"),
   311 => (x"b2",x"73",x"33",x"c2"),
   312 => (x"97",x"e8",x"da",x"c2"),
   313 => (x"c0",x"c3",x"4b",x"bf"),
   314 => (x"2b",x"b7",x"c6",x"9b"),
   315 => (x"81",x"c2",x"b2",x"73"),
   316 => (x"30",x"71",x"48",x"c1"),
   317 => (x"48",x"c1",x"49",x"70"),
   318 => (x"4d",x"70",x"30",x"75"),
   319 => (x"84",x"c1",x"4c",x"72"),
   320 => (x"c0",x"c8",x"94",x"71"),
   321 => (x"cc",x"06",x"ad",x"b7"),
   322 => (x"b7",x"34",x"c1",x"87"),
   323 => (x"b7",x"c0",x"c8",x"2d"),
   324 => (x"f4",x"ff",x"01",x"ad"),
   325 => (x"f0",x"48",x"74",x"87"),
   326 => (x"5e",x"0e",x"87",x"d7"),
   327 => (x"0e",x"5d",x"5c",x"5b"),
   328 => (x"e3",x"c2",x"86",x"f8"),
   329 => (x"78",x"c0",x"48",x"c6"),
   330 => (x"1e",x"fe",x"da",x"c2"),
   331 => (x"de",x"fb",x"49",x"c0"),
   332 => (x"70",x"86",x"c4",x"87"),
   333 => (x"87",x"c5",x"05",x"98"),
   334 => (x"c0",x"c9",x"48",x"c0"),
   335 => (x"c1",x"4d",x"c0",x"87"),
   336 => (x"dd",x"f2",x"c0",x"7e"),
   337 => (x"db",x"c2",x"49",x"bf"),
   338 => (x"c8",x"71",x"4a",x"f4"),
   339 => (x"87",x"d9",x"ec",x"4b"),
   340 => (x"c2",x"05",x"98",x"70"),
   341 => (x"c0",x"7e",x"c0",x"87"),
   342 => (x"49",x"bf",x"d9",x"f2"),
   343 => (x"4a",x"d0",x"dc",x"c2"),
   344 => (x"ec",x"4b",x"c8",x"71"),
   345 => (x"98",x"70",x"87",x"c3"),
   346 => (x"c0",x"87",x"c2",x"05"),
   347 => (x"c0",x"02",x"6e",x"7e"),
   348 => (x"e2",x"c2",x"87",x"fd"),
   349 => (x"c2",x"4d",x"bf",x"c4"),
   350 => (x"bf",x"9f",x"fc",x"e2"),
   351 => (x"d6",x"c5",x"48",x"7e"),
   352 => (x"c7",x"05",x"a8",x"ea"),
   353 => (x"c4",x"e2",x"c2",x"87"),
   354 => (x"87",x"ce",x"4d",x"bf"),
   355 => (x"e9",x"ca",x"48",x"6e"),
   356 => (x"c5",x"02",x"a8",x"d5"),
   357 => (x"c7",x"48",x"c0",x"87"),
   358 => (x"da",x"c2",x"87",x"e3"),
   359 => (x"49",x"75",x"1e",x"fe"),
   360 => (x"c4",x"87",x"ec",x"f9"),
   361 => (x"05",x"98",x"70",x"86"),
   362 => (x"48",x"c0",x"87",x"c5"),
   363 => (x"c0",x"87",x"ce",x"c7"),
   364 => (x"49",x"bf",x"d9",x"f2"),
   365 => (x"4a",x"d0",x"dc",x"c2"),
   366 => (x"ea",x"4b",x"c8",x"71"),
   367 => (x"98",x"70",x"87",x"eb"),
   368 => (x"c2",x"87",x"c8",x"05"),
   369 => (x"c1",x"48",x"c6",x"e3"),
   370 => (x"c0",x"87",x"da",x"78"),
   371 => (x"49",x"bf",x"dd",x"f2"),
   372 => (x"4a",x"f4",x"db",x"c2"),
   373 => (x"ea",x"4b",x"c8",x"71"),
   374 => (x"98",x"70",x"87",x"cf"),
   375 => (x"87",x"c5",x"c0",x"02"),
   376 => (x"d8",x"c6",x"48",x"c0"),
   377 => (x"fc",x"e2",x"c2",x"87"),
   378 => (x"c1",x"49",x"bf",x"97"),
   379 => (x"c0",x"05",x"a9",x"d5"),
   380 => (x"e2",x"c2",x"87",x"cd"),
   381 => (x"49",x"bf",x"97",x"fd"),
   382 => (x"02",x"a9",x"ea",x"c2"),
   383 => (x"c0",x"87",x"c5",x"c0"),
   384 => (x"87",x"f9",x"c5",x"48"),
   385 => (x"97",x"fe",x"da",x"c2"),
   386 => (x"c3",x"48",x"7e",x"bf"),
   387 => (x"c0",x"02",x"a8",x"e9"),
   388 => (x"48",x"6e",x"87",x"ce"),
   389 => (x"02",x"a8",x"eb",x"c3"),
   390 => (x"c0",x"87",x"c5",x"c0"),
   391 => (x"87",x"dd",x"c5",x"48"),
   392 => (x"97",x"c9",x"db",x"c2"),
   393 => (x"05",x"99",x"49",x"bf"),
   394 => (x"c2",x"87",x"cc",x"c0"),
   395 => (x"bf",x"97",x"ca",x"db"),
   396 => (x"02",x"a9",x"c2",x"49"),
   397 => (x"c0",x"87",x"c5",x"c0"),
   398 => (x"87",x"c1",x"c5",x"48"),
   399 => (x"97",x"cb",x"db",x"c2"),
   400 => (x"e3",x"c2",x"48",x"bf"),
   401 => (x"4c",x"70",x"58",x"c2"),
   402 => (x"c2",x"88",x"c1",x"48"),
   403 => (x"c2",x"58",x"c6",x"e3"),
   404 => (x"bf",x"97",x"cc",x"db"),
   405 => (x"c2",x"81",x"75",x"49"),
   406 => (x"bf",x"97",x"cd",x"db"),
   407 => (x"72",x"32",x"c8",x"4a"),
   408 => (x"e7",x"c2",x"7e",x"a1"),
   409 => (x"78",x"6e",x"48",x"d3"),
   410 => (x"97",x"ce",x"db",x"c2"),
   411 => (x"a6",x"c8",x"48",x"bf"),
   412 => (x"c6",x"e3",x"c2",x"58"),
   413 => (x"cf",x"c2",x"02",x"bf"),
   414 => (x"d9",x"f2",x"c0",x"87"),
   415 => (x"dc",x"c2",x"49",x"bf"),
   416 => (x"c8",x"71",x"4a",x"d0"),
   417 => (x"87",x"e1",x"e7",x"4b"),
   418 => (x"c0",x"02",x"98",x"70"),
   419 => (x"48",x"c0",x"87",x"c5"),
   420 => (x"c2",x"87",x"ea",x"c3"),
   421 => (x"4c",x"bf",x"fe",x"e2"),
   422 => (x"5c",x"e7",x"e7",x"c2"),
   423 => (x"97",x"e3",x"db",x"c2"),
   424 => (x"31",x"c8",x"49",x"bf"),
   425 => (x"97",x"e2",x"db",x"c2"),
   426 => (x"49",x"a1",x"4a",x"bf"),
   427 => (x"97",x"e4",x"db",x"c2"),
   428 => (x"32",x"d0",x"4a",x"bf"),
   429 => (x"c2",x"49",x"a1",x"72"),
   430 => (x"bf",x"97",x"e5",x"db"),
   431 => (x"72",x"32",x"d8",x"4a"),
   432 => (x"66",x"c4",x"49",x"a1"),
   433 => (x"d3",x"e7",x"c2",x"91"),
   434 => (x"e7",x"c2",x"81",x"bf"),
   435 => (x"db",x"c2",x"59",x"db"),
   436 => (x"4a",x"bf",x"97",x"eb"),
   437 => (x"db",x"c2",x"32",x"c8"),
   438 => (x"4b",x"bf",x"97",x"ea"),
   439 => (x"db",x"c2",x"4a",x"a2"),
   440 => (x"4b",x"bf",x"97",x"ec"),
   441 => (x"a2",x"73",x"33",x"d0"),
   442 => (x"ed",x"db",x"c2",x"4a"),
   443 => (x"cf",x"4b",x"bf",x"97"),
   444 => (x"73",x"33",x"d8",x"9b"),
   445 => (x"e7",x"c2",x"4a",x"a2"),
   446 => (x"8a",x"c2",x"5a",x"df"),
   447 => (x"e7",x"c2",x"92",x"74"),
   448 => (x"a1",x"72",x"48",x"df"),
   449 => (x"87",x"c1",x"c1",x"78"),
   450 => (x"97",x"d0",x"db",x"c2"),
   451 => (x"31",x"c8",x"49",x"bf"),
   452 => (x"97",x"cf",x"db",x"c2"),
   453 => (x"49",x"a1",x"4a",x"bf"),
   454 => (x"ff",x"c7",x"31",x"c5"),
   455 => (x"c2",x"29",x"c9",x"81"),
   456 => (x"c2",x"59",x"e7",x"e7"),
   457 => (x"bf",x"97",x"d5",x"db"),
   458 => (x"c2",x"32",x"c8",x"4a"),
   459 => (x"bf",x"97",x"d4",x"db"),
   460 => (x"c4",x"4a",x"a2",x"4b"),
   461 => (x"82",x"6e",x"92",x"66"),
   462 => (x"5a",x"e3",x"e7",x"c2"),
   463 => (x"48",x"db",x"e7",x"c2"),
   464 => (x"e7",x"c2",x"78",x"c0"),
   465 => (x"a1",x"72",x"48",x"d7"),
   466 => (x"e7",x"e7",x"c2",x"78"),
   467 => (x"db",x"e7",x"c2",x"48"),
   468 => (x"e7",x"c2",x"78",x"bf"),
   469 => (x"e7",x"c2",x"48",x"eb"),
   470 => (x"c2",x"78",x"bf",x"df"),
   471 => (x"02",x"bf",x"c6",x"e3"),
   472 => (x"74",x"87",x"c9",x"c0"),
   473 => (x"70",x"30",x"c4",x"48"),
   474 => (x"87",x"c9",x"c0",x"7e"),
   475 => (x"bf",x"e3",x"e7",x"c2"),
   476 => (x"70",x"30",x"c4",x"48"),
   477 => (x"ca",x"e3",x"c2",x"7e"),
   478 => (x"c1",x"78",x"6e",x"48"),
   479 => (x"26",x"8e",x"f8",x"48"),
   480 => (x"26",x"4c",x"26",x"4d"),
   481 => (x"0e",x"4f",x"26",x"4b"),
   482 => (x"5d",x"5c",x"5b",x"5e"),
   483 => (x"c2",x"4a",x"71",x"0e"),
   484 => (x"02",x"bf",x"c6",x"e3"),
   485 => (x"4b",x"72",x"87",x"cb"),
   486 => (x"4d",x"72",x"2b",x"c7"),
   487 => (x"c9",x"9d",x"ff",x"c1"),
   488 => (x"c8",x"4b",x"72",x"87"),
   489 => (x"c3",x"4d",x"72",x"2b"),
   490 => (x"e7",x"c2",x"9d",x"ff"),
   491 => (x"c0",x"83",x"bf",x"d3"),
   492 => (x"ab",x"bf",x"d5",x"f2"),
   493 => (x"c0",x"87",x"d9",x"02"),
   494 => (x"c2",x"5b",x"d9",x"f2"),
   495 => (x"73",x"1e",x"fe",x"da"),
   496 => (x"87",x"cb",x"f1",x"49"),
   497 => (x"98",x"70",x"86",x"c4"),
   498 => (x"c0",x"87",x"c5",x"05"),
   499 => (x"87",x"e6",x"c0",x"48"),
   500 => (x"bf",x"c6",x"e3",x"c2"),
   501 => (x"75",x"87",x"d2",x"02"),
   502 => (x"c2",x"91",x"c4",x"49"),
   503 => (x"69",x"81",x"fe",x"da"),
   504 => (x"ff",x"ff",x"cf",x"4c"),
   505 => (x"cb",x"9c",x"ff",x"ff"),
   506 => (x"c2",x"49",x"75",x"87"),
   507 => (x"fe",x"da",x"c2",x"91"),
   508 => (x"4c",x"69",x"9f",x"81"),
   509 => (x"c6",x"fe",x"48",x"74"),
   510 => (x"5b",x"5e",x"0e",x"87"),
   511 => (x"f8",x"0e",x"5d",x"5c"),
   512 => (x"9c",x"4c",x"71",x"86"),
   513 => (x"c0",x"87",x"c5",x"05"),
   514 => (x"87",x"c0",x"c3",x"48"),
   515 => (x"48",x"7e",x"a4",x"c8"),
   516 => (x"66",x"d8",x"78",x"c0"),
   517 => (x"d8",x"87",x"c7",x"02"),
   518 => (x"05",x"bf",x"97",x"66"),
   519 => (x"48",x"c0",x"87",x"c5"),
   520 => (x"c0",x"87",x"e9",x"c2"),
   521 => (x"49",x"49",x"c1",x"1e"),
   522 => (x"c4",x"87",x"d3",x"ca"),
   523 => (x"9d",x"4d",x"70",x"86"),
   524 => (x"87",x"c2",x"c1",x"02"),
   525 => (x"4a",x"ce",x"e3",x"c2"),
   526 => (x"e0",x"49",x"66",x"d8"),
   527 => (x"98",x"70",x"87",x"d0"),
   528 => (x"87",x"f2",x"c0",x"02"),
   529 => (x"66",x"d8",x"4a",x"75"),
   530 => (x"e0",x"4b",x"cb",x"49"),
   531 => (x"98",x"70",x"87",x"f5"),
   532 => (x"87",x"e2",x"c0",x"02"),
   533 => (x"9d",x"75",x"1e",x"c0"),
   534 => (x"c8",x"87",x"c7",x"02"),
   535 => (x"78",x"c0",x"48",x"a6"),
   536 => (x"a6",x"c8",x"87",x"c5"),
   537 => (x"c8",x"78",x"c1",x"48"),
   538 => (x"d1",x"c9",x"49",x"66"),
   539 => (x"70",x"86",x"c4",x"87"),
   540 => (x"fe",x"05",x"9d",x"4d"),
   541 => (x"9d",x"75",x"87",x"fe"),
   542 => (x"87",x"ce",x"c1",x"02"),
   543 => (x"6e",x"49",x"a5",x"dc"),
   544 => (x"da",x"78",x"69",x"48"),
   545 => (x"a6",x"c4",x"49",x"a5"),
   546 => (x"78",x"a4",x"c4",x"48"),
   547 => (x"c4",x"48",x"69",x"9f"),
   548 => (x"c2",x"78",x"08",x"66"),
   549 => (x"02",x"bf",x"c6",x"e3"),
   550 => (x"a5",x"d4",x"87",x"d2"),
   551 => (x"49",x"69",x"9f",x"49"),
   552 => (x"99",x"ff",x"ff",x"c0"),
   553 => (x"30",x"d0",x"48",x"71"),
   554 => (x"87",x"c2",x"7e",x"70"),
   555 => (x"48",x"6e",x"7e",x"c0"),
   556 => (x"80",x"bf",x"66",x"c4"),
   557 => (x"78",x"08",x"66",x"c4"),
   558 => (x"a4",x"cc",x"7c",x"c0"),
   559 => (x"bf",x"66",x"c4",x"49"),
   560 => (x"49",x"a4",x"d0",x"79"),
   561 => (x"48",x"c1",x"79",x"c0"),
   562 => (x"48",x"c0",x"87",x"c2"),
   563 => (x"ee",x"fa",x"8e",x"f8"),
   564 => (x"5b",x"5e",x"0e",x"87"),
   565 => (x"4c",x"71",x"0e",x"5c"),
   566 => (x"cb",x"c1",x"02",x"9c"),
   567 => (x"49",x"a4",x"c8",x"87"),
   568 => (x"c3",x"c1",x"02",x"69"),
   569 => (x"cc",x"49",x"6c",x"87"),
   570 => (x"80",x"71",x"48",x"66"),
   571 => (x"70",x"58",x"a6",x"d0"),
   572 => (x"c2",x"e3",x"c2",x"b9"),
   573 => (x"ba",x"ff",x"4a",x"bf"),
   574 => (x"99",x"71",x"99",x"72"),
   575 => (x"87",x"e5",x"c0",x"02"),
   576 => (x"6b",x"4b",x"a4",x"c4"),
   577 => (x"87",x"ff",x"f9",x"49"),
   578 => (x"e2",x"c2",x"7b",x"70"),
   579 => (x"6c",x"49",x"bf",x"fe"),
   580 => (x"cc",x"7c",x"71",x"81"),
   581 => (x"e3",x"c2",x"b9",x"66"),
   582 => (x"ff",x"4a",x"bf",x"c2"),
   583 => (x"71",x"99",x"72",x"ba"),
   584 => (x"db",x"ff",x"05",x"99"),
   585 => (x"7c",x"66",x"cc",x"87"),
   586 => (x"1e",x"87",x"d6",x"f9"),
   587 => (x"4b",x"71",x"1e",x"73"),
   588 => (x"87",x"c7",x"02",x"9b"),
   589 => (x"69",x"49",x"a3",x"c8"),
   590 => (x"c0",x"87",x"c5",x"05"),
   591 => (x"87",x"f6",x"c0",x"48"),
   592 => (x"bf",x"d7",x"e7",x"c2"),
   593 => (x"4a",x"a3",x"c4",x"49"),
   594 => (x"8a",x"c2",x"4a",x"6a"),
   595 => (x"bf",x"fe",x"e2",x"c2"),
   596 => (x"49",x"a1",x"72",x"92"),
   597 => (x"bf",x"c2",x"e3",x"c2"),
   598 => (x"72",x"9a",x"6b",x"4a"),
   599 => (x"f2",x"c0",x"49",x"a1"),
   600 => (x"66",x"c8",x"59",x"d9"),
   601 => (x"e6",x"ea",x"71",x"1e"),
   602 => (x"70",x"86",x"c4",x"87"),
   603 => (x"87",x"c4",x"05",x"98"),
   604 => (x"87",x"c2",x"48",x"c0"),
   605 => (x"ca",x"f8",x"48",x"c1"),
   606 => (x"1e",x"73",x"1e",x"87"),
   607 => (x"02",x"9b",x"4b",x"71"),
   608 => (x"a3",x"c8",x"87",x"c7"),
   609 => (x"c5",x"05",x"69",x"49"),
   610 => (x"c0",x"48",x"c0",x"87"),
   611 => (x"e7",x"c2",x"87",x"f6"),
   612 => (x"c4",x"49",x"bf",x"d7"),
   613 => (x"4a",x"6a",x"4a",x"a3"),
   614 => (x"e2",x"c2",x"8a",x"c2"),
   615 => (x"72",x"92",x"bf",x"fe"),
   616 => (x"e3",x"c2",x"49",x"a1"),
   617 => (x"6b",x"4a",x"bf",x"c2"),
   618 => (x"49",x"a1",x"72",x"9a"),
   619 => (x"59",x"d9",x"f2",x"c0"),
   620 => (x"71",x"1e",x"66",x"c8"),
   621 => (x"c4",x"87",x"d1",x"e6"),
   622 => (x"05",x"98",x"70",x"86"),
   623 => (x"48",x"c0",x"87",x"c4"),
   624 => (x"48",x"c1",x"87",x"c2"),
   625 => (x"0e",x"87",x"fc",x"f6"),
   626 => (x"5d",x"5c",x"5b",x"5e"),
   627 => (x"4b",x"71",x"1e",x"0e"),
   628 => (x"73",x"4d",x"66",x"d4"),
   629 => (x"cc",x"c1",x"02",x"9b"),
   630 => (x"49",x"a3",x"c8",x"87"),
   631 => (x"c4",x"c1",x"02",x"69"),
   632 => (x"4c",x"a3",x"d0",x"87"),
   633 => (x"bf",x"c2",x"e3",x"c2"),
   634 => (x"6c",x"b9",x"ff",x"49"),
   635 => (x"d4",x"7e",x"99",x"4a"),
   636 => (x"cd",x"06",x"a9",x"66"),
   637 => (x"7c",x"7b",x"c0",x"87"),
   638 => (x"c4",x"4a",x"a3",x"cc"),
   639 => (x"79",x"6a",x"49",x"a3"),
   640 => (x"49",x"72",x"87",x"ca"),
   641 => (x"d4",x"99",x"c0",x"f8"),
   642 => (x"8d",x"71",x"4d",x"66"),
   643 => (x"29",x"c9",x"49",x"75"),
   644 => (x"49",x"73",x"1e",x"71"),
   645 => (x"c2",x"87",x"fa",x"fa"),
   646 => (x"73",x"1e",x"fe",x"da"),
   647 => (x"87",x"cb",x"fc",x"49"),
   648 => (x"66",x"d4",x"86",x"c8"),
   649 => (x"d6",x"f5",x"26",x"7c"),
   650 => (x"1e",x"73",x"1e",x"87"),
   651 => (x"02",x"9b",x"4b",x"71"),
   652 => (x"c2",x"87",x"e4",x"c0"),
   653 => (x"73",x"5b",x"eb",x"e7"),
   654 => (x"c2",x"8a",x"c2",x"4a"),
   655 => (x"49",x"bf",x"fe",x"e2"),
   656 => (x"d7",x"e7",x"c2",x"92"),
   657 => (x"80",x"72",x"48",x"bf"),
   658 => (x"58",x"ef",x"e7",x"c2"),
   659 => (x"30",x"c4",x"48",x"71"),
   660 => (x"58",x"ce",x"e3",x"c2"),
   661 => (x"c2",x"87",x"ed",x"c0"),
   662 => (x"c2",x"48",x"e7",x"e7"),
   663 => (x"78",x"bf",x"db",x"e7"),
   664 => (x"48",x"eb",x"e7",x"c2"),
   665 => (x"bf",x"df",x"e7",x"c2"),
   666 => (x"c6",x"e3",x"c2",x"78"),
   667 => (x"87",x"c9",x"02",x"bf"),
   668 => (x"bf",x"fe",x"e2",x"c2"),
   669 => (x"c7",x"31",x"c4",x"49"),
   670 => (x"e3",x"e7",x"c2",x"87"),
   671 => (x"31",x"c4",x"49",x"bf"),
   672 => (x"59",x"ce",x"e3",x"c2"),
   673 => (x"0e",x"87",x"fc",x"f3"),
   674 => (x"0e",x"5c",x"5b",x"5e"),
   675 => (x"4b",x"c0",x"4a",x"71"),
   676 => (x"c0",x"02",x"9a",x"72"),
   677 => (x"a2",x"da",x"87",x"e0"),
   678 => (x"4b",x"69",x"9f",x"49"),
   679 => (x"bf",x"c6",x"e3",x"c2"),
   680 => (x"d4",x"87",x"cf",x"02"),
   681 => (x"69",x"9f",x"49",x"a2"),
   682 => (x"ff",x"c0",x"4c",x"49"),
   683 => (x"34",x"d0",x"9c",x"ff"),
   684 => (x"4c",x"c0",x"87",x"c2"),
   685 => (x"49",x"73",x"b3",x"74"),
   686 => (x"f3",x"87",x"ee",x"fd"),
   687 => (x"5e",x"0e",x"87",x"c3"),
   688 => (x"0e",x"5d",x"5c",x"5b"),
   689 => (x"4a",x"71",x"86",x"f4"),
   690 => (x"9a",x"72",x"7e",x"c0"),
   691 => (x"c2",x"87",x"d8",x"02"),
   692 => (x"c0",x"48",x"fa",x"da"),
   693 => (x"f2",x"da",x"c2",x"78"),
   694 => (x"eb",x"e7",x"c2",x"48"),
   695 => (x"da",x"c2",x"78",x"bf"),
   696 => (x"e7",x"c2",x"48",x"f6"),
   697 => (x"c2",x"78",x"bf",x"e7"),
   698 => (x"c0",x"48",x"db",x"e3"),
   699 => (x"ca",x"e3",x"c2",x"50"),
   700 => (x"da",x"c2",x"49",x"bf"),
   701 => (x"71",x"4a",x"bf",x"fa"),
   702 => (x"c9",x"c4",x"03",x"aa"),
   703 => (x"cf",x"49",x"72",x"87"),
   704 => (x"e9",x"c0",x"05",x"99"),
   705 => (x"d5",x"f2",x"c0",x"87"),
   706 => (x"f2",x"da",x"c2",x"48"),
   707 => (x"da",x"c2",x"78",x"bf"),
   708 => (x"da",x"c2",x"1e",x"fe"),
   709 => (x"c2",x"49",x"bf",x"f2"),
   710 => (x"c1",x"48",x"f2",x"da"),
   711 => (x"e3",x"71",x"78",x"a1"),
   712 => (x"86",x"c4",x"87",x"ed"),
   713 => (x"48",x"d1",x"f2",x"c0"),
   714 => (x"78",x"fe",x"da",x"c2"),
   715 => (x"f2",x"c0",x"87",x"cc"),
   716 => (x"c0",x"48",x"bf",x"d1"),
   717 => (x"f2",x"c0",x"80",x"e0"),
   718 => (x"da",x"c2",x"58",x"d5"),
   719 => (x"c1",x"48",x"bf",x"fa"),
   720 => (x"fe",x"da",x"c2",x"80"),
   721 => (x"0c",x"91",x"27",x"58"),
   722 => (x"97",x"bf",x"00",x"00"),
   723 => (x"02",x"9d",x"4d",x"bf"),
   724 => (x"c3",x"87",x"e3",x"c2"),
   725 => (x"c2",x"02",x"ad",x"e5"),
   726 => (x"f2",x"c0",x"87",x"dc"),
   727 => (x"cb",x"4b",x"bf",x"d1"),
   728 => (x"4c",x"11",x"49",x"a3"),
   729 => (x"c1",x"05",x"ac",x"cf"),
   730 => (x"49",x"75",x"87",x"d2"),
   731 => (x"89",x"c1",x"99",x"df"),
   732 => (x"e3",x"c2",x"91",x"cd"),
   733 => (x"a3",x"c1",x"81",x"ce"),
   734 => (x"c3",x"51",x"12",x"4a"),
   735 => (x"51",x"12",x"4a",x"a3"),
   736 => (x"12",x"4a",x"a3",x"c5"),
   737 => (x"4a",x"a3",x"c7",x"51"),
   738 => (x"a3",x"c9",x"51",x"12"),
   739 => (x"ce",x"51",x"12",x"4a"),
   740 => (x"51",x"12",x"4a",x"a3"),
   741 => (x"12",x"4a",x"a3",x"d0"),
   742 => (x"4a",x"a3",x"d2",x"51"),
   743 => (x"a3",x"d4",x"51",x"12"),
   744 => (x"d6",x"51",x"12",x"4a"),
   745 => (x"51",x"12",x"4a",x"a3"),
   746 => (x"12",x"4a",x"a3",x"d8"),
   747 => (x"4a",x"a3",x"dc",x"51"),
   748 => (x"a3",x"de",x"51",x"12"),
   749 => (x"c1",x"51",x"12",x"4a"),
   750 => (x"87",x"fa",x"c0",x"7e"),
   751 => (x"99",x"c8",x"49",x"74"),
   752 => (x"87",x"eb",x"c0",x"05"),
   753 => (x"99",x"d0",x"49",x"74"),
   754 => (x"dc",x"87",x"d1",x"05"),
   755 => (x"cb",x"c0",x"02",x"66"),
   756 => (x"dc",x"49",x"73",x"87"),
   757 => (x"98",x"70",x"0f",x"66"),
   758 => (x"87",x"d3",x"c0",x"02"),
   759 => (x"c6",x"c0",x"05",x"6e"),
   760 => (x"ce",x"e3",x"c2",x"87"),
   761 => (x"c0",x"50",x"c0",x"48"),
   762 => (x"48",x"bf",x"d1",x"f2"),
   763 => (x"c2",x"87",x"dd",x"c2"),
   764 => (x"c0",x"48",x"db",x"e3"),
   765 => (x"e3",x"c2",x"7e",x"50"),
   766 => (x"c2",x"49",x"bf",x"ca"),
   767 => (x"4a",x"bf",x"fa",x"da"),
   768 => (x"fb",x"04",x"aa",x"71"),
   769 => (x"e7",x"c2",x"87",x"f7"),
   770 => (x"c0",x"05",x"bf",x"eb"),
   771 => (x"e3",x"c2",x"87",x"c8"),
   772 => (x"c1",x"02",x"bf",x"c6"),
   773 => (x"da",x"c2",x"87",x"f4"),
   774 => (x"ed",x"49",x"bf",x"f6"),
   775 => (x"da",x"c2",x"87",x"e9"),
   776 => (x"a6",x"c4",x"58",x"fa"),
   777 => (x"f6",x"da",x"c2",x"48"),
   778 => (x"e3",x"c2",x"78",x"bf"),
   779 => (x"c0",x"02",x"bf",x"c6"),
   780 => (x"66",x"c4",x"87",x"d8"),
   781 => (x"ff",x"ff",x"cf",x"49"),
   782 => (x"a9",x"99",x"f8",x"ff"),
   783 => (x"87",x"c5",x"c0",x"02"),
   784 => (x"e1",x"c0",x"4c",x"c0"),
   785 => (x"c0",x"4c",x"c1",x"87"),
   786 => (x"66",x"c4",x"87",x"dc"),
   787 => (x"f8",x"ff",x"cf",x"49"),
   788 => (x"c0",x"02",x"a9",x"99"),
   789 => (x"a6",x"c8",x"87",x"c8"),
   790 => (x"c0",x"78",x"c0",x"48"),
   791 => (x"a6",x"c8",x"87",x"c5"),
   792 => (x"c8",x"78",x"c1",x"48"),
   793 => (x"9c",x"74",x"4c",x"66"),
   794 => (x"87",x"de",x"c0",x"05"),
   795 => (x"c2",x"49",x"66",x"c4"),
   796 => (x"fe",x"e2",x"c2",x"89"),
   797 => (x"e7",x"c2",x"91",x"bf"),
   798 => (x"71",x"48",x"bf",x"d7"),
   799 => (x"f6",x"da",x"c2",x"80"),
   800 => (x"fa",x"da",x"c2",x"58"),
   801 => (x"f9",x"78",x"c0",x"48"),
   802 => (x"48",x"c0",x"87",x"e3"),
   803 => (x"ee",x"eb",x"8e",x"f4"),
   804 => (x"00",x"00",x"00",x"87"),
   805 => (x"ff",x"ff",x"ff",x"00"),
   806 => (x"00",x"0c",x"a1",x"ff"),
   807 => (x"00",x"0c",x"aa",x"00"),
   808 => (x"54",x"41",x"46",x"00"),
   809 => (x"20",x"20",x"32",x"33"),
   810 => (x"41",x"46",x"00",x"20"),
   811 => (x"20",x"36",x"31",x"54"),
   812 => (x"1e",x"00",x"20",x"20"),
   813 => (x"c3",x"48",x"d4",x"ff"),
   814 => (x"48",x"68",x"78",x"ff"),
   815 => (x"ff",x"1e",x"4f",x"26"),
   816 => (x"ff",x"c3",x"48",x"d4"),
   817 => (x"48",x"d0",x"ff",x"78"),
   818 => (x"ff",x"78",x"e1",x"c0"),
   819 => (x"78",x"d4",x"48",x"d4"),
   820 => (x"48",x"ef",x"e7",x"c2"),
   821 => (x"50",x"bf",x"d4",x"ff"),
   822 => (x"ff",x"1e",x"4f",x"26"),
   823 => (x"e0",x"c0",x"48",x"d0"),
   824 => (x"1e",x"4f",x"26",x"78"),
   825 => (x"70",x"87",x"cc",x"ff"),
   826 => (x"c6",x"02",x"99",x"49"),
   827 => (x"a9",x"fb",x"c0",x"87"),
   828 => (x"71",x"87",x"f1",x"05"),
   829 => (x"0e",x"4f",x"26",x"48"),
   830 => (x"0e",x"5c",x"5b",x"5e"),
   831 => (x"4c",x"c0",x"4b",x"71"),
   832 => (x"70",x"87",x"f0",x"fe"),
   833 => (x"c0",x"02",x"99",x"49"),
   834 => (x"ec",x"c0",x"87",x"f9"),
   835 => (x"f2",x"c0",x"02",x"a9"),
   836 => (x"a9",x"fb",x"c0",x"87"),
   837 => (x"87",x"eb",x"c0",x"02"),
   838 => (x"ac",x"b7",x"66",x"cc"),
   839 => (x"d0",x"87",x"c7",x"03"),
   840 => (x"87",x"c2",x"02",x"66"),
   841 => (x"99",x"71",x"53",x"71"),
   842 => (x"c1",x"87",x"c2",x"02"),
   843 => (x"87",x"c3",x"fe",x"84"),
   844 => (x"02",x"99",x"49",x"70"),
   845 => (x"ec",x"c0",x"87",x"cd"),
   846 => (x"87",x"c7",x"02",x"a9"),
   847 => (x"05",x"a9",x"fb",x"c0"),
   848 => (x"d0",x"87",x"d5",x"ff"),
   849 => (x"87",x"c3",x"02",x"66"),
   850 => (x"c0",x"7b",x"97",x"c0"),
   851 => (x"c4",x"05",x"a9",x"ec"),
   852 => (x"c5",x"4a",x"74",x"87"),
   853 => (x"c0",x"4a",x"74",x"87"),
   854 => (x"48",x"72",x"8a",x"0a"),
   855 => (x"4d",x"26",x"87",x"c2"),
   856 => (x"4b",x"26",x"4c",x"26"),
   857 => (x"fd",x"1e",x"4f",x"26"),
   858 => (x"4a",x"70",x"87",x"c9"),
   859 => (x"04",x"aa",x"f0",x"c0"),
   860 => (x"f9",x"c0",x"87",x"c9"),
   861 => (x"87",x"c3",x"01",x"aa"),
   862 => (x"c1",x"8a",x"f0",x"c0"),
   863 => (x"c9",x"04",x"aa",x"c1"),
   864 => (x"aa",x"da",x"c1",x"87"),
   865 => (x"c0",x"87",x"c3",x"01"),
   866 => (x"48",x"72",x"8a",x"f7"),
   867 => (x"5e",x"0e",x"4f",x"26"),
   868 => (x"71",x"0e",x"5c",x"5b"),
   869 => (x"4b",x"d4",x"ff",x"4a"),
   870 => (x"e7",x"c0",x"49",x"72"),
   871 => (x"9c",x"4c",x"70",x"87"),
   872 => (x"c1",x"87",x"c2",x"02"),
   873 => (x"48",x"d0",x"ff",x"8c"),
   874 => (x"d5",x"c1",x"78",x"c5"),
   875 => (x"c6",x"49",x"74",x"7b"),
   876 => (x"ee",x"e3",x"c1",x"31"),
   877 => (x"48",x"4a",x"bf",x"97"),
   878 => (x"7b",x"70",x"b0",x"71"),
   879 => (x"c4",x"48",x"d0",x"ff"),
   880 => (x"87",x"dc",x"fe",x"78"),
   881 => (x"5c",x"5b",x"5e",x"0e"),
   882 => (x"86",x"f8",x"0e",x"5d"),
   883 => (x"7e",x"c0",x"4c",x"71"),
   884 => (x"c0",x"87",x"eb",x"fb"),
   885 => (x"f1",x"f9",x"c0",x"4b"),
   886 => (x"c0",x"49",x"bf",x"97"),
   887 => (x"87",x"cf",x"04",x"a9"),
   888 => (x"c1",x"87",x"c0",x"fc"),
   889 => (x"f1",x"f9",x"c0",x"83"),
   890 => (x"ab",x"49",x"bf",x"97"),
   891 => (x"c0",x"87",x"f1",x"06"),
   892 => (x"bf",x"97",x"f1",x"f9"),
   893 => (x"fa",x"87",x"cf",x"02"),
   894 => (x"49",x"70",x"87",x"f9"),
   895 => (x"87",x"c6",x"02",x"99"),
   896 => (x"05",x"a9",x"ec",x"c0"),
   897 => (x"4b",x"c0",x"87",x"f1"),
   898 => (x"70",x"87",x"e8",x"fa"),
   899 => (x"87",x"e3",x"fa",x"4d"),
   900 => (x"fa",x"58",x"a6",x"c8"),
   901 => (x"4a",x"70",x"87",x"dd"),
   902 => (x"a4",x"c8",x"83",x"c1"),
   903 => (x"49",x"69",x"97",x"49"),
   904 => (x"87",x"c7",x"02",x"ad"),
   905 => (x"05",x"ad",x"ff",x"c0"),
   906 => (x"c9",x"87",x"e7",x"c0"),
   907 => (x"69",x"97",x"49",x"a4"),
   908 => (x"a9",x"66",x"c4",x"49"),
   909 => (x"48",x"87",x"c7",x"02"),
   910 => (x"05",x"a8",x"ff",x"c0"),
   911 => (x"a4",x"ca",x"87",x"d4"),
   912 => (x"49",x"69",x"97",x"49"),
   913 => (x"87",x"c6",x"02",x"aa"),
   914 => (x"05",x"aa",x"ff",x"c0"),
   915 => (x"7e",x"c1",x"87",x"c4"),
   916 => (x"ec",x"c0",x"87",x"d0"),
   917 => (x"87",x"c6",x"02",x"ad"),
   918 => (x"05",x"ad",x"fb",x"c0"),
   919 => (x"4b",x"c0",x"87",x"c4"),
   920 => (x"02",x"6e",x"7e",x"c1"),
   921 => (x"f9",x"87",x"e1",x"fe"),
   922 => (x"48",x"73",x"87",x"f0"),
   923 => (x"ed",x"fb",x"8e",x"f8"),
   924 => (x"5e",x"0e",x"00",x"87"),
   925 => (x"0e",x"5d",x"5c",x"5b"),
   926 => (x"4d",x"71",x"86",x"f8"),
   927 => (x"75",x"4b",x"d4",x"ff"),
   928 => (x"f4",x"e7",x"c2",x"1e"),
   929 => (x"87",x"f1",x"e5",x"49"),
   930 => (x"98",x"70",x"86",x"c4"),
   931 => (x"87",x"ca",x"c4",x"02"),
   932 => (x"c1",x"48",x"a6",x"c4"),
   933 => (x"78",x"bf",x"f0",x"e3"),
   934 => (x"f1",x"fb",x"49",x"75"),
   935 => (x"48",x"d0",x"ff",x"87"),
   936 => (x"d6",x"c1",x"78",x"c5"),
   937 => (x"75",x"4a",x"c0",x"7b"),
   938 => (x"7b",x"11",x"49",x"a2"),
   939 => (x"b7",x"cb",x"82",x"c1"),
   940 => (x"87",x"f3",x"04",x"aa"),
   941 => (x"ff",x"c3",x"4a",x"cc"),
   942 => (x"c0",x"82",x"c1",x"7b"),
   943 => (x"04",x"aa",x"b7",x"e0"),
   944 => (x"d0",x"ff",x"87",x"f4"),
   945 => (x"c3",x"78",x"c4",x"48"),
   946 => (x"78",x"c5",x"7b",x"ff"),
   947 => (x"c1",x"7b",x"d3",x"c1"),
   948 => (x"66",x"78",x"c4",x"7b"),
   949 => (x"a8",x"b7",x"c0",x"48"),
   950 => (x"87",x"ee",x"c2",x"06"),
   951 => (x"bf",x"fc",x"e7",x"c2"),
   952 => (x"48",x"66",x"c4",x"4c"),
   953 => (x"a6",x"c8",x"88",x"74"),
   954 => (x"02",x"9c",x"74",x"58"),
   955 => (x"c2",x"87",x"f7",x"c1"),
   956 => (x"c8",x"7e",x"fe",x"da"),
   957 => (x"c0",x"8c",x"4d",x"c0"),
   958 => (x"c6",x"03",x"ac",x"b7"),
   959 => (x"a4",x"c0",x"c8",x"87"),
   960 => (x"c2",x"4c",x"c0",x"4d"),
   961 => (x"bf",x"97",x"ef",x"e7"),
   962 => (x"02",x"99",x"d0",x"49"),
   963 => (x"1e",x"c0",x"87",x"d0"),
   964 => (x"49",x"f4",x"e7",x"c2"),
   965 => (x"c4",x"87",x"d4",x"e8"),
   966 => (x"c0",x"4a",x"70",x"86"),
   967 => (x"da",x"c2",x"87",x"ed"),
   968 => (x"e7",x"c2",x"1e",x"fe"),
   969 => (x"c2",x"e8",x"49",x"f4"),
   970 => (x"70",x"86",x"c4",x"87"),
   971 => (x"48",x"d0",x"ff",x"4a"),
   972 => (x"c1",x"78",x"c5",x"c8"),
   973 => (x"97",x"6e",x"7b",x"d4"),
   974 => (x"48",x"6e",x"7b",x"bf"),
   975 => (x"7e",x"70",x"80",x"c1"),
   976 => (x"ff",x"05",x"8d",x"c1"),
   977 => (x"d0",x"ff",x"87",x"f0"),
   978 => (x"72",x"78",x"c4",x"48"),
   979 => (x"87",x"c5",x"05",x"9a"),
   980 => (x"c7",x"c1",x"48",x"c0"),
   981 => (x"c2",x"1e",x"c1",x"87"),
   982 => (x"e5",x"49",x"f4",x"e7"),
   983 => (x"86",x"c4",x"87",x"f3"),
   984 => (x"fe",x"05",x"9c",x"74"),
   985 => (x"66",x"c4",x"87",x"c9"),
   986 => (x"a8",x"b7",x"c0",x"48"),
   987 => (x"c2",x"87",x"d1",x"06"),
   988 => (x"c0",x"48",x"f4",x"e7"),
   989 => (x"c0",x"80",x"d0",x"78"),
   990 => (x"c2",x"80",x"f4",x"78"),
   991 => (x"78",x"bf",x"c0",x"e8"),
   992 => (x"c0",x"48",x"66",x"c4"),
   993 => (x"fd",x"01",x"a8",x"b7"),
   994 => (x"d0",x"ff",x"87",x"d2"),
   995 => (x"c1",x"78",x"c5",x"48"),
   996 => (x"7b",x"c0",x"7b",x"d3"),
   997 => (x"48",x"c1",x"78",x"c4"),
   998 => (x"48",x"c0",x"87",x"c2"),
   999 => (x"4d",x"26",x"8e",x"f8"),
  1000 => (x"4b",x"26",x"4c",x"26"),
  1001 => (x"5e",x"0e",x"4f",x"26"),
  1002 => (x"0e",x"5d",x"5c",x"5b"),
  1003 => (x"c0",x"4b",x"71",x"1e"),
  1004 => (x"04",x"ab",x"4d",x"4c"),
  1005 => (x"c0",x"87",x"e8",x"c0"),
  1006 => (x"75",x"1e",x"c4",x"f7"),
  1007 => (x"87",x"c4",x"02",x"9d"),
  1008 => (x"87",x"c2",x"4a",x"c0"),
  1009 => (x"49",x"72",x"4a",x"c1"),
  1010 => (x"c4",x"87",x"f3",x"eb"),
  1011 => (x"c1",x"7e",x"70",x"86"),
  1012 => (x"c2",x"05",x"6e",x"84"),
  1013 => (x"c1",x"4c",x"73",x"87"),
  1014 => (x"06",x"ac",x"73",x"85"),
  1015 => (x"6e",x"87",x"d8",x"ff"),
  1016 => (x"f9",x"fe",x"26",x"48"),
  1017 => (x"5b",x"5e",x"0e",x"87"),
  1018 => (x"4b",x"71",x"0e",x"5c"),
  1019 => (x"d8",x"02",x"66",x"cc"),
  1020 => (x"f0",x"c0",x"4c",x"87"),
  1021 => (x"87",x"d8",x"02",x"8c"),
  1022 => (x"8a",x"c1",x"4a",x"74"),
  1023 => (x"8a",x"87",x"d1",x"02"),
  1024 => (x"8a",x"87",x"cd",x"02"),
  1025 => (x"d9",x"87",x"c9",x"02"),
  1026 => (x"f9",x"49",x"73",x"87"),
  1027 => (x"87",x"d2",x"87",x"e4"),
  1028 => (x"49",x"c0",x"1e",x"74"),
  1029 => (x"87",x"f5",x"d7",x"c1"),
  1030 => (x"49",x"73",x"1e",x"74"),
  1031 => (x"87",x"ed",x"d7",x"c1"),
  1032 => (x"fb",x"fd",x"86",x"c8"),
  1033 => (x"5b",x"5e",x"0e",x"87"),
  1034 => (x"1e",x"0e",x"5d",x"5c"),
  1035 => (x"de",x"49",x"4c",x"71"),
  1036 => (x"dc",x"e8",x"c2",x"91"),
  1037 => (x"97",x"85",x"71",x"4d"),
  1038 => (x"dc",x"c1",x"02",x"6d"),
  1039 => (x"c8",x"e8",x"c2",x"87"),
  1040 => (x"81",x"74",x"49",x"bf"),
  1041 => (x"87",x"de",x"fd",x"71"),
  1042 => (x"98",x"48",x"7e",x"70"),
  1043 => (x"87",x"f2",x"c0",x"02"),
  1044 => (x"4b",x"d0",x"e8",x"c2"),
  1045 => (x"49",x"cb",x"4a",x"70"),
  1046 => (x"87",x"cb",x"c1",x"ff"),
  1047 => (x"93",x"cb",x"4b",x"74"),
  1048 => (x"83",x"c2",x"e4",x"c1"),
  1049 => (x"c2",x"c1",x"83",x"c4"),
  1050 => (x"49",x"74",x"7b",x"dd"),
  1051 => (x"87",x"cb",x"c1",x"c1"),
  1052 => (x"e3",x"c1",x"7b",x"75"),
  1053 => (x"49",x"bf",x"97",x"ef"),
  1054 => (x"d0",x"e8",x"c2",x"1e"),
  1055 => (x"87",x"e5",x"fd",x"49"),
  1056 => (x"49",x"74",x"86",x"c4"),
  1057 => (x"87",x"f3",x"c0",x"c1"),
  1058 => (x"c2",x"c1",x"49",x"c0"),
  1059 => (x"e7",x"c2",x"87",x"d2"),
  1060 => (x"78",x"c0",x"48",x"f0"),
  1061 => (x"fb",x"dd",x"49",x"c1"),
  1062 => (x"c1",x"fc",x"26",x"87"),
  1063 => (x"61",x"6f",x"4c",x"87"),
  1064 => (x"67",x"6e",x"69",x"64"),
  1065 => (x"00",x"2e",x"2e",x"2e"),
  1066 => (x"71",x"1e",x"73",x"1e"),
  1067 => (x"e8",x"c2",x"49",x"4a"),
  1068 => (x"71",x"81",x"bf",x"c8"),
  1069 => (x"70",x"87",x"ef",x"fb"),
  1070 => (x"c4",x"02",x"9b",x"4b"),
  1071 => (x"c6",x"e7",x"49",x"87"),
  1072 => (x"c8",x"e8",x"c2",x"87"),
  1073 => (x"c1",x"78",x"c0",x"48"),
  1074 => (x"87",x"c8",x"dd",x"49"),
  1075 => (x"1e",x"87",x"d3",x"fb"),
  1076 => (x"c1",x"c1",x"49",x"c0"),
  1077 => (x"4f",x"26",x"87",x"ca"),
  1078 => (x"49",x"4a",x"71",x"1e"),
  1079 => (x"e4",x"c1",x"91",x"cb"),
  1080 => (x"81",x"c8",x"81",x"c2"),
  1081 => (x"e7",x"c2",x"48",x"11"),
  1082 => (x"e8",x"c2",x"58",x"f4"),
  1083 => (x"78",x"c0",x"48",x"c8"),
  1084 => (x"df",x"dc",x"49",x"c1"),
  1085 => (x"1e",x"4f",x"26",x"87"),
  1086 => (x"d2",x"02",x"99",x"71"),
  1087 => (x"d7",x"e5",x"c1",x"87"),
  1088 => (x"f7",x"50",x"c0",x"48"),
  1089 => (x"d8",x"c3",x"c1",x"80"),
  1090 => (x"fb",x"e3",x"c1",x"40"),
  1091 => (x"c1",x"87",x"ce",x"78"),
  1092 => (x"c1",x"48",x"d3",x"e5"),
  1093 => (x"fc",x"78",x"f4",x"e3"),
  1094 => (x"cf",x"c3",x"c1",x"80"),
  1095 => (x"0e",x"4f",x"26",x"78"),
  1096 => (x"5d",x"5c",x"5b",x"5e"),
  1097 => (x"c2",x"86",x"f4",x"0e"),
  1098 => (x"c0",x"4d",x"fe",x"da"),
  1099 => (x"48",x"a6",x"c4",x"4c"),
  1100 => (x"e8",x"c2",x"78",x"c0"),
  1101 => (x"c0",x"48",x"bf",x"c8"),
  1102 => (x"c0",x"c1",x"06",x"a8"),
  1103 => (x"fe",x"da",x"c2",x"87"),
  1104 => (x"c0",x"02",x"98",x"48"),
  1105 => (x"f7",x"c0",x"87",x"f7"),
  1106 => (x"66",x"c8",x"1e",x"c4"),
  1107 => (x"c4",x"87",x"c7",x"02"),
  1108 => (x"78",x"c0",x"48",x"a6"),
  1109 => (x"a6",x"c4",x"87",x"c5"),
  1110 => (x"c4",x"78",x"c1",x"48"),
  1111 => (x"dd",x"e5",x"49",x"66"),
  1112 => (x"70",x"86",x"c4",x"87"),
  1113 => (x"c4",x"84",x"c1",x"4d"),
  1114 => (x"80",x"c1",x"48",x"66"),
  1115 => (x"c2",x"58",x"a6",x"c8"),
  1116 => (x"ac",x"bf",x"c8",x"e8"),
  1117 => (x"75",x"87",x"c6",x"03"),
  1118 => (x"c9",x"ff",x"05",x"9d"),
  1119 => (x"75",x"4c",x"c0",x"87"),
  1120 => (x"dc",x"c3",x"02",x"9d"),
  1121 => (x"c4",x"f7",x"c0",x"87"),
  1122 => (x"02",x"66",x"c8",x"1e"),
  1123 => (x"a6",x"cc",x"87",x"c7"),
  1124 => (x"c5",x"78",x"c0",x"48"),
  1125 => (x"48",x"a6",x"cc",x"87"),
  1126 => (x"66",x"cc",x"78",x"c1"),
  1127 => (x"87",x"de",x"e4",x"49"),
  1128 => (x"7e",x"70",x"86",x"c4"),
  1129 => (x"c2",x"02",x"98",x"48"),
  1130 => (x"cb",x"49",x"87",x"e4"),
  1131 => (x"49",x"69",x"97",x"81"),
  1132 => (x"c1",x"02",x"99",x"d0"),
  1133 => (x"49",x"74",x"87",x"d4"),
  1134 => (x"e4",x"c1",x"91",x"cb"),
  1135 => (x"c2",x"c1",x"81",x"c2"),
  1136 => (x"81",x"c8",x"79",x"e8"),
  1137 => (x"74",x"51",x"ff",x"c3"),
  1138 => (x"c2",x"91",x"de",x"49"),
  1139 => (x"71",x"4d",x"dc",x"e8"),
  1140 => (x"97",x"c1",x"c2",x"85"),
  1141 => (x"49",x"a5",x"c1",x"7d"),
  1142 => (x"c2",x"51",x"e0",x"c0"),
  1143 => (x"bf",x"97",x"ce",x"e3"),
  1144 => (x"c1",x"87",x"d2",x"02"),
  1145 => (x"4b",x"a5",x"c2",x"84"),
  1146 => (x"4a",x"ce",x"e3",x"c2"),
  1147 => (x"fa",x"fe",x"49",x"db"),
  1148 => (x"d9",x"c1",x"87",x"f5"),
  1149 => (x"49",x"a5",x"cd",x"87"),
  1150 => (x"84",x"c1",x"51",x"c0"),
  1151 => (x"6e",x"4b",x"a5",x"c2"),
  1152 => (x"fe",x"49",x"cb",x"4a"),
  1153 => (x"c1",x"87",x"e0",x"fa"),
  1154 => (x"49",x"74",x"87",x"c4"),
  1155 => (x"e4",x"c1",x"91",x"cb"),
  1156 => (x"c0",x"c1",x"81",x"c2"),
  1157 => (x"e3",x"c2",x"79",x"e5"),
  1158 => (x"02",x"bf",x"97",x"ce"),
  1159 => (x"49",x"74",x"87",x"d8"),
  1160 => (x"84",x"c1",x"91",x"de"),
  1161 => (x"4b",x"dc",x"e8",x"c2"),
  1162 => (x"e3",x"c2",x"83",x"71"),
  1163 => (x"49",x"dd",x"4a",x"ce"),
  1164 => (x"87",x"f3",x"f9",x"fe"),
  1165 => (x"4b",x"74",x"87",x"d8"),
  1166 => (x"e8",x"c2",x"93",x"de"),
  1167 => (x"a3",x"cb",x"83",x"dc"),
  1168 => (x"c1",x"51",x"c0",x"49"),
  1169 => (x"4a",x"6e",x"73",x"84"),
  1170 => (x"f9",x"fe",x"49",x"cb"),
  1171 => (x"66",x"c4",x"87",x"d9"),
  1172 => (x"c8",x"80",x"c1",x"48"),
  1173 => (x"ac",x"c7",x"58",x"a6"),
  1174 => (x"87",x"c5",x"c0",x"03"),
  1175 => (x"e4",x"fc",x"05",x"6e"),
  1176 => (x"f4",x"48",x"74",x"87"),
  1177 => (x"87",x"f6",x"f4",x"8e"),
  1178 => (x"71",x"1e",x"73",x"1e"),
  1179 => (x"91",x"cb",x"49",x"4b"),
  1180 => (x"81",x"c2",x"e4",x"c1"),
  1181 => (x"c1",x"4a",x"a1",x"c8"),
  1182 => (x"12",x"48",x"ee",x"e3"),
  1183 => (x"4a",x"a1",x"c9",x"50"),
  1184 => (x"48",x"f1",x"f9",x"c0"),
  1185 => (x"81",x"ca",x"50",x"12"),
  1186 => (x"48",x"ef",x"e3",x"c1"),
  1187 => (x"e3",x"c1",x"50",x"11"),
  1188 => (x"49",x"bf",x"97",x"ef"),
  1189 => (x"f5",x"49",x"c0",x"1e"),
  1190 => (x"e7",x"c2",x"87",x"cb"),
  1191 => (x"78",x"de",x"48",x"f0"),
  1192 => (x"ef",x"d5",x"49",x"c1"),
  1193 => (x"f9",x"f3",x"26",x"87"),
  1194 => (x"5b",x"5e",x"0e",x"87"),
  1195 => (x"f4",x"0e",x"5d",x"5c"),
  1196 => (x"49",x"4d",x"71",x"86"),
  1197 => (x"e4",x"c1",x"91",x"cb"),
  1198 => (x"a1",x"c8",x"81",x"c2"),
  1199 => (x"7e",x"a1",x"ca",x"4a"),
  1200 => (x"c2",x"48",x"a6",x"c4"),
  1201 => (x"78",x"bf",x"f8",x"eb"),
  1202 => (x"4b",x"bf",x"97",x"6e"),
  1203 => (x"73",x"4c",x"66",x"c4"),
  1204 => (x"cc",x"48",x"12",x"2c"),
  1205 => (x"9c",x"70",x"58",x"a6"),
  1206 => (x"81",x"c9",x"84",x"c1"),
  1207 => (x"b7",x"49",x"69",x"97"),
  1208 => (x"87",x"c2",x"04",x"ac"),
  1209 => (x"97",x"6e",x"4c",x"c0"),
  1210 => (x"66",x"c8",x"4a",x"bf"),
  1211 => (x"ff",x"31",x"72",x"49"),
  1212 => (x"99",x"66",x"c4",x"b9"),
  1213 => (x"30",x"72",x"48",x"74"),
  1214 => (x"71",x"48",x"4a",x"70"),
  1215 => (x"fc",x"eb",x"c2",x"b0"),
  1216 => (x"f6",x"e4",x"c0",x"58"),
  1217 => (x"d4",x"49",x"c0",x"87"),
  1218 => (x"49",x"75",x"87",x"ca"),
  1219 => (x"87",x"eb",x"f6",x"c0"),
  1220 => (x"c9",x"f2",x"8e",x"f4"),
  1221 => (x"1e",x"73",x"1e",x"87"),
  1222 => (x"fe",x"49",x"4b",x"71"),
  1223 => (x"49",x"73",x"87",x"cb"),
  1224 => (x"f1",x"87",x"c6",x"fe"),
  1225 => (x"73",x"1e",x"87",x"fc"),
  1226 => (x"c6",x"4b",x"71",x"1e"),
  1227 => (x"db",x"02",x"4a",x"a3"),
  1228 => (x"02",x"8a",x"c1",x"87"),
  1229 => (x"02",x"8a",x"87",x"d6"),
  1230 => (x"8a",x"87",x"da",x"c1"),
  1231 => (x"87",x"fc",x"c0",x"02"),
  1232 => (x"e1",x"c0",x"02",x"8a"),
  1233 => (x"cb",x"02",x"8a",x"87"),
  1234 => (x"87",x"db",x"c1",x"87"),
  1235 => (x"c7",x"f6",x"49",x"c7"),
  1236 => (x"87",x"de",x"c1",x"87"),
  1237 => (x"bf",x"c8",x"e8",x"c2"),
  1238 => (x"87",x"cb",x"c1",x"02"),
  1239 => (x"c2",x"88",x"c1",x"48"),
  1240 => (x"c1",x"58",x"cc",x"e8"),
  1241 => (x"e8",x"c2",x"87",x"c1"),
  1242 => (x"c0",x"02",x"bf",x"cc"),
  1243 => (x"e8",x"c2",x"87",x"f9"),
  1244 => (x"c1",x"48",x"bf",x"c8"),
  1245 => (x"cc",x"e8",x"c2",x"80"),
  1246 => (x"87",x"eb",x"c0",x"58"),
  1247 => (x"bf",x"c8",x"e8",x"c2"),
  1248 => (x"c2",x"89",x"c6",x"49"),
  1249 => (x"c0",x"59",x"cc",x"e8"),
  1250 => (x"da",x"03",x"a9",x"b7"),
  1251 => (x"c8",x"e8",x"c2",x"87"),
  1252 => (x"d2",x"78",x"c0",x"48"),
  1253 => (x"cc",x"e8",x"c2",x"87"),
  1254 => (x"87",x"cb",x"02",x"bf"),
  1255 => (x"bf",x"c8",x"e8",x"c2"),
  1256 => (x"c2",x"80",x"c6",x"48"),
  1257 => (x"c0",x"58",x"cc",x"e8"),
  1258 => (x"87",x"e8",x"d1",x"49"),
  1259 => (x"f4",x"c0",x"49",x"73"),
  1260 => (x"ed",x"ef",x"87",x"c9"),
  1261 => (x"5b",x"5e",x"0e",x"87"),
  1262 => (x"ff",x"0e",x"5d",x"5c"),
  1263 => (x"a6",x"dc",x"86",x"d4"),
  1264 => (x"48",x"a6",x"c8",x"59"),
  1265 => (x"80",x"c4",x"78",x"c0"),
  1266 => (x"78",x"66",x"c0",x"c1"),
  1267 => (x"78",x"c1",x"80",x"c4"),
  1268 => (x"78",x"c1",x"80",x"c4"),
  1269 => (x"48",x"cc",x"e8",x"c2"),
  1270 => (x"e7",x"c2",x"78",x"c1"),
  1271 => (x"de",x"48",x"bf",x"f0"),
  1272 => (x"87",x"c9",x"05",x"a8"),
  1273 => (x"cc",x"87",x"f8",x"f4"),
  1274 => (x"e6",x"cf",x"58",x"a6"),
  1275 => (x"87",x"ce",x"e3",x"87"),
  1276 => (x"e2",x"87",x"f0",x"e3"),
  1277 => (x"4c",x"70",x"87",x"fd"),
  1278 => (x"02",x"ac",x"fb",x"c0"),
  1279 => (x"d8",x"87",x"fb",x"c1"),
  1280 => (x"ed",x"c1",x"05",x"66"),
  1281 => (x"66",x"fc",x"c0",x"87"),
  1282 => (x"6a",x"82",x"c4",x"4a"),
  1283 => (x"c1",x"1e",x"72",x"7e"),
  1284 => (x"c4",x"48",x"c8",x"e0"),
  1285 => (x"a1",x"c8",x"49",x"66"),
  1286 => (x"71",x"41",x"20",x"4a"),
  1287 => (x"87",x"f9",x"05",x"aa"),
  1288 => (x"4a",x"26",x"51",x"10"),
  1289 => (x"48",x"66",x"fc",x"c0"),
  1290 => (x"78",x"e8",x"c9",x"c1"),
  1291 => (x"81",x"c7",x"49",x"6a"),
  1292 => (x"fc",x"c0",x"51",x"74"),
  1293 => (x"81",x"c8",x"49",x"66"),
  1294 => (x"fc",x"c0",x"51",x"c1"),
  1295 => (x"81",x"c9",x"49",x"66"),
  1296 => (x"fc",x"c0",x"51",x"c0"),
  1297 => (x"81",x"ca",x"49",x"66"),
  1298 => (x"1e",x"c1",x"51",x"c0"),
  1299 => (x"49",x"6a",x"1e",x"d8"),
  1300 => (x"e2",x"e2",x"81",x"c8"),
  1301 => (x"c1",x"86",x"c8",x"87"),
  1302 => (x"c0",x"48",x"66",x"c0"),
  1303 => (x"87",x"c7",x"01",x"a8"),
  1304 => (x"c1",x"48",x"a6",x"c8"),
  1305 => (x"c1",x"87",x"ce",x"78"),
  1306 => (x"c1",x"48",x"66",x"c0"),
  1307 => (x"58",x"a6",x"d0",x"88"),
  1308 => (x"ee",x"e1",x"87",x"c3"),
  1309 => (x"48",x"a6",x"d0",x"87"),
  1310 => (x"9c",x"74",x"78",x"c2"),
  1311 => (x"87",x"cf",x"cd",x"02"),
  1312 => (x"c1",x"48",x"66",x"c8"),
  1313 => (x"03",x"a8",x"66",x"c4"),
  1314 => (x"dc",x"87",x"c4",x"cd"),
  1315 => (x"78",x"c0",x"48",x"a6"),
  1316 => (x"78",x"c0",x"80",x"e8"),
  1317 => (x"70",x"87",x"dc",x"e0"),
  1318 => (x"ac",x"d0",x"c1",x"4c"),
  1319 => (x"87",x"d7",x"c2",x"05"),
  1320 => (x"e3",x"7e",x"66",x"c4"),
  1321 => (x"a6",x"c8",x"87",x"c0"),
  1322 => (x"87",x"c7",x"e0",x"58"),
  1323 => (x"ec",x"c0",x"4c",x"70"),
  1324 => (x"ed",x"c1",x"05",x"ac"),
  1325 => (x"49",x"66",x"c8",x"87"),
  1326 => (x"fc",x"c0",x"91",x"cb"),
  1327 => (x"a1",x"c4",x"81",x"66"),
  1328 => (x"c8",x"4d",x"6a",x"4a"),
  1329 => (x"66",x"c4",x"4a",x"a1"),
  1330 => (x"d8",x"c3",x"c1",x"52"),
  1331 => (x"e2",x"df",x"ff",x"79"),
  1332 => (x"9c",x"4c",x"70",x"87"),
  1333 => (x"c0",x"87",x"d9",x"02"),
  1334 => (x"d3",x"02",x"ac",x"fb"),
  1335 => (x"ff",x"55",x"74",x"87"),
  1336 => (x"70",x"87",x"d0",x"df"),
  1337 => (x"c7",x"02",x"9c",x"4c"),
  1338 => (x"ac",x"fb",x"c0",x"87"),
  1339 => (x"87",x"ed",x"ff",x"05"),
  1340 => (x"c2",x"55",x"e0",x"c0"),
  1341 => (x"97",x"c0",x"55",x"c1"),
  1342 => (x"48",x"66",x"d8",x"7d"),
  1343 => (x"db",x"05",x"a8",x"6e"),
  1344 => (x"48",x"66",x"c8",x"87"),
  1345 => (x"04",x"a8",x"66",x"cc"),
  1346 => (x"66",x"c8",x"87",x"ca"),
  1347 => (x"cc",x"80",x"c1",x"48"),
  1348 => (x"87",x"c8",x"58",x"a6"),
  1349 => (x"c1",x"48",x"66",x"cc"),
  1350 => (x"58",x"a6",x"d0",x"88"),
  1351 => (x"87",x"d3",x"de",x"ff"),
  1352 => (x"d0",x"c1",x"4c",x"70"),
  1353 => (x"87",x"c8",x"05",x"ac"),
  1354 => (x"c1",x"48",x"66",x"d4"),
  1355 => (x"58",x"a6",x"d8",x"80"),
  1356 => (x"02",x"ac",x"d0",x"c1"),
  1357 => (x"c4",x"87",x"e9",x"fd"),
  1358 => (x"66",x"d8",x"48",x"66"),
  1359 => (x"e0",x"c9",x"05",x"a8"),
  1360 => (x"a6",x"e0",x"c0",x"87"),
  1361 => (x"74",x"78",x"c0",x"48"),
  1362 => (x"88",x"fb",x"c0",x"48"),
  1363 => (x"98",x"48",x"7e",x"70"),
  1364 => (x"87",x"e2",x"c9",x"02"),
  1365 => (x"70",x"88",x"cb",x"48"),
  1366 => (x"02",x"98",x"48",x"7e"),
  1367 => (x"48",x"87",x"cd",x"c1"),
  1368 => (x"7e",x"70",x"88",x"c9"),
  1369 => (x"c3",x"02",x"98",x"48"),
  1370 => (x"c4",x"48",x"87",x"fe"),
  1371 => (x"48",x"7e",x"70",x"88"),
  1372 => (x"87",x"ce",x"02",x"98"),
  1373 => (x"70",x"88",x"c1",x"48"),
  1374 => (x"02",x"98",x"48",x"7e"),
  1375 => (x"c8",x"87",x"e9",x"c3"),
  1376 => (x"a6",x"dc",x"87",x"d6"),
  1377 => (x"78",x"f0",x"c0",x"48"),
  1378 => (x"87",x"e7",x"dc",x"ff"),
  1379 => (x"ec",x"c0",x"4c",x"70"),
  1380 => (x"c4",x"c0",x"02",x"ac"),
  1381 => (x"a6",x"e0",x"c0",x"87"),
  1382 => (x"ac",x"ec",x"c0",x"5c"),
  1383 => (x"ff",x"87",x"cd",x"02"),
  1384 => (x"70",x"87",x"d0",x"dc"),
  1385 => (x"ac",x"ec",x"c0",x"4c"),
  1386 => (x"87",x"f3",x"ff",x"05"),
  1387 => (x"02",x"ac",x"ec",x"c0"),
  1388 => (x"ff",x"87",x"c4",x"c0"),
  1389 => (x"c0",x"87",x"fc",x"db"),
  1390 => (x"d0",x"1e",x"ca",x"1e"),
  1391 => (x"91",x"cb",x"49",x"66"),
  1392 => (x"48",x"66",x"c4",x"c1"),
  1393 => (x"a6",x"cc",x"80",x"71"),
  1394 => (x"48",x"66",x"c8",x"58"),
  1395 => (x"a6",x"d0",x"80",x"c4"),
  1396 => (x"bf",x"66",x"cc",x"58"),
  1397 => (x"de",x"dc",x"ff",x"49"),
  1398 => (x"de",x"1e",x"c1",x"87"),
  1399 => (x"bf",x"66",x"d4",x"1e"),
  1400 => (x"d2",x"dc",x"ff",x"49"),
  1401 => (x"70",x"86",x"d0",x"87"),
  1402 => (x"08",x"c0",x"48",x"49"),
  1403 => (x"a6",x"e8",x"c0",x"88"),
  1404 => (x"06",x"a8",x"c0",x"58"),
  1405 => (x"c0",x"87",x"ee",x"c0"),
  1406 => (x"dd",x"48",x"66",x"e4"),
  1407 => (x"e4",x"c0",x"03",x"a8"),
  1408 => (x"bf",x"66",x"c4",x"87"),
  1409 => (x"66",x"e4",x"c0",x"49"),
  1410 => (x"51",x"e0",x"c0",x"81"),
  1411 => (x"49",x"66",x"e4",x"c0"),
  1412 => (x"66",x"c4",x"81",x"c1"),
  1413 => (x"c1",x"c2",x"81",x"bf"),
  1414 => (x"66",x"e4",x"c0",x"51"),
  1415 => (x"c4",x"81",x"c2",x"49"),
  1416 => (x"c0",x"81",x"bf",x"66"),
  1417 => (x"c1",x"48",x"6e",x"51"),
  1418 => (x"6e",x"78",x"e8",x"c9"),
  1419 => (x"d0",x"81",x"c8",x"49"),
  1420 => (x"49",x"6e",x"51",x"66"),
  1421 => (x"66",x"d4",x"81",x"c9"),
  1422 => (x"ca",x"49",x"6e",x"51"),
  1423 => (x"51",x"66",x"dc",x"81"),
  1424 => (x"c1",x"48",x"66",x"d0"),
  1425 => (x"58",x"a6",x"d4",x"80"),
  1426 => (x"cc",x"48",x"66",x"c8"),
  1427 => (x"c0",x"04",x"a8",x"66"),
  1428 => (x"66",x"c8",x"87",x"cb"),
  1429 => (x"cc",x"80",x"c1",x"48"),
  1430 => (x"d9",x"c5",x"58",x"a6"),
  1431 => (x"48",x"66",x"cc",x"87"),
  1432 => (x"a6",x"d0",x"88",x"c1"),
  1433 => (x"87",x"ce",x"c5",x"58"),
  1434 => (x"87",x"fa",x"db",x"ff"),
  1435 => (x"58",x"a6",x"e8",x"c0"),
  1436 => (x"87",x"f2",x"db",x"ff"),
  1437 => (x"58",x"a6",x"e0",x"c0"),
  1438 => (x"05",x"a8",x"ec",x"c0"),
  1439 => (x"dc",x"87",x"ca",x"c0"),
  1440 => (x"e4",x"c0",x"48",x"a6"),
  1441 => (x"c4",x"c0",x"78",x"66"),
  1442 => (x"e6",x"d8",x"ff",x"87"),
  1443 => (x"49",x"66",x"c8",x"87"),
  1444 => (x"fc",x"c0",x"91",x"cb"),
  1445 => (x"80",x"71",x"48",x"66"),
  1446 => (x"c8",x"4a",x"7e",x"70"),
  1447 => (x"ca",x"49",x"6e",x"82"),
  1448 => (x"66",x"e4",x"c0",x"81"),
  1449 => (x"49",x"66",x"dc",x"51"),
  1450 => (x"e4",x"c0",x"81",x"c1"),
  1451 => (x"48",x"c1",x"89",x"66"),
  1452 => (x"49",x"70",x"30",x"71"),
  1453 => (x"97",x"71",x"89",x"c1"),
  1454 => (x"f8",x"eb",x"c2",x"7a"),
  1455 => (x"e4",x"c0",x"49",x"bf"),
  1456 => (x"6a",x"97",x"29",x"66"),
  1457 => (x"98",x"71",x"48",x"4a"),
  1458 => (x"58",x"a6",x"ec",x"c0"),
  1459 => (x"81",x"c4",x"49",x"6e"),
  1460 => (x"66",x"d8",x"4d",x"69"),
  1461 => (x"a8",x"66",x"c4",x"48"),
  1462 => (x"87",x"c8",x"c0",x"02"),
  1463 => (x"c0",x"48",x"a6",x"c4"),
  1464 => (x"87",x"c5",x"c0",x"78"),
  1465 => (x"c1",x"48",x"a6",x"c4"),
  1466 => (x"1e",x"66",x"c4",x"78"),
  1467 => (x"75",x"1e",x"e0",x"c0"),
  1468 => (x"c2",x"d8",x"ff",x"49"),
  1469 => (x"70",x"86",x"c8",x"87"),
  1470 => (x"ac",x"b7",x"c0",x"4c"),
  1471 => (x"87",x"d4",x"c1",x"06"),
  1472 => (x"e0",x"c0",x"85",x"74"),
  1473 => (x"75",x"89",x"74",x"49"),
  1474 => (x"d1",x"e0",x"c1",x"4b"),
  1475 => (x"e6",x"fe",x"71",x"4a"),
  1476 => (x"85",x"c2",x"87",x"d5"),
  1477 => (x"48",x"66",x"e0",x"c0"),
  1478 => (x"e4",x"c0",x"80",x"c1"),
  1479 => (x"e8",x"c0",x"58",x"a6"),
  1480 => (x"81",x"c1",x"49",x"66"),
  1481 => (x"c0",x"02",x"a9",x"70"),
  1482 => (x"a6",x"c4",x"87",x"c8"),
  1483 => (x"c0",x"78",x"c0",x"48"),
  1484 => (x"a6",x"c4",x"87",x"c5"),
  1485 => (x"c4",x"78",x"c1",x"48"),
  1486 => (x"a4",x"c2",x"1e",x"66"),
  1487 => (x"48",x"e0",x"c0",x"49"),
  1488 => (x"49",x"70",x"88",x"71"),
  1489 => (x"ff",x"49",x"75",x"1e"),
  1490 => (x"c8",x"87",x"ec",x"d6"),
  1491 => (x"a8",x"b7",x"c0",x"86"),
  1492 => (x"87",x"c0",x"ff",x"01"),
  1493 => (x"02",x"66",x"e0",x"c0"),
  1494 => (x"6e",x"87",x"d1",x"c0"),
  1495 => (x"c0",x"81",x"c9",x"49"),
  1496 => (x"6e",x"51",x"66",x"e0"),
  1497 => (x"e9",x"ca",x"c1",x"48"),
  1498 => (x"87",x"cc",x"c0",x"78"),
  1499 => (x"81",x"c9",x"49",x"6e"),
  1500 => (x"48",x"6e",x"51",x"c2"),
  1501 => (x"78",x"d5",x"cc",x"c1"),
  1502 => (x"cc",x"48",x"66",x"c8"),
  1503 => (x"c0",x"04",x"a8",x"66"),
  1504 => (x"66",x"c8",x"87",x"cb"),
  1505 => (x"cc",x"80",x"c1",x"48"),
  1506 => (x"e9",x"c0",x"58",x"a6"),
  1507 => (x"48",x"66",x"cc",x"87"),
  1508 => (x"a6",x"d0",x"88",x"c1"),
  1509 => (x"87",x"de",x"c0",x"58"),
  1510 => (x"87",x"c7",x"d5",x"ff"),
  1511 => (x"d5",x"c0",x"4c",x"70"),
  1512 => (x"ac",x"c6",x"c1",x"87"),
  1513 => (x"87",x"c8",x"c0",x"05"),
  1514 => (x"c1",x"48",x"66",x"d0"),
  1515 => (x"58",x"a6",x"d4",x"80"),
  1516 => (x"87",x"ef",x"d4",x"ff"),
  1517 => (x"66",x"d4",x"4c",x"70"),
  1518 => (x"d8",x"80",x"c1",x"48"),
  1519 => (x"9c",x"74",x"58",x"a6"),
  1520 => (x"87",x"cb",x"c0",x"02"),
  1521 => (x"c1",x"48",x"66",x"c8"),
  1522 => (x"04",x"a8",x"66",x"c4"),
  1523 => (x"ff",x"87",x"fc",x"f2"),
  1524 => (x"c8",x"87",x"c7",x"d4"),
  1525 => (x"a8",x"c7",x"48",x"66"),
  1526 => (x"87",x"e5",x"c0",x"03"),
  1527 => (x"48",x"cc",x"e8",x"c2"),
  1528 => (x"66",x"c8",x"78",x"c0"),
  1529 => (x"c0",x"91",x"cb",x"49"),
  1530 => (x"c4",x"81",x"66",x"fc"),
  1531 => (x"4a",x"6a",x"4a",x"a1"),
  1532 => (x"c8",x"79",x"52",x"c0"),
  1533 => (x"80",x"c1",x"48",x"66"),
  1534 => (x"c7",x"58",x"a6",x"cc"),
  1535 => (x"db",x"ff",x"04",x"a8"),
  1536 => (x"8e",x"d4",x"ff",x"87"),
  1537 => (x"87",x"d6",x"de",x"ff"),
  1538 => (x"64",x"61",x"6f",x"4c"),
  1539 => (x"20",x"2e",x"2a",x"20"),
  1540 => (x"00",x"20",x"3a",x"00"),
  1541 => (x"71",x"1e",x"73",x"1e"),
  1542 => (x"c6",x"02",x"9b",x"4b"),
  1543 => (x"c8",x"e8",x"c2",x"87"),
  1544 => (x"c7",x"78",x"c0",x"48"),
  1545 => (x"c8",x"e8",x"c2",x"1e"),
  1546 => (x"e4",x"c1",x"1e",x"bf"),
  1547 => (x"e7",x"c2",x"1e",x"c2"),
  1548 => (x"ed",x"49",x"bf",x"f0"),
  1549 => (x"86",x"cc",x"87",x"ff"),
  1550 => (x"bf",x"f0",x"e7",x"c2"),
  1551 => (x"87",x"f7",x"e2",x"49"),
  1552 => (x"c8",x"02",x"9b",x"73"),
  1553 => (x"c2",x"e4",x"c1",x"87"),
  1554 => (x"c0",x"e3",x"c0",x"49"),
  1555 => (x"d1",x"dd",x"ff",x"87"),
  1556 => (x"e3",x"c1",x"1e",x"87"),
  1557 => (x"50",x"c0",x"48",x"ee"),
  1558 => (x"bf",x"e5",x"e5",x"c1"),
  1559 => (x"d1",x"d8",x"ff",x"49"),
  1560 => (x"26",x"48",x"c0",x"87"),
  1561 => (x"e3",x"c7",x"1e",x"4f"),
  1562 => (x"fe",x"49",x"c1",x"87"),
  1563 => (x"e9",x"fe",x"87",x"e6"),
  1564 => (x"98",x"70",x"87",x"e5"),
  1565 => (x"fe",x"87",x"cd",x"02"),
  1566 => (x"70",x"87",x"df",x"f2"),
  1567 => (x"87",x"c4",x"02",x"98"),
  1568 => (x"87",x"c2",x"4a",x"c1"),
  1569 => (x"9a",x"72",x"4a",x"c0"),
  1570 => (x"c0",x"87",x"ce",x"05"),
  1571 => (x"f5",x"e2",x"c1",x"1e"),
  1572 => (x"ee",x"ee",x"c0",x"49"),
  1573 => (x"fe",x"86",x"c4",x"87"),
  1574 => (x"c1",x"1e",x"c0",x"87"),
  1575 => (x"c0",x"49",x"c0",x"e3"),
  1576 => (x"c0",x"87",x"e0",x"ee"),
  1577 => (x"87",x"e9",x"fe",x"1e"),
  1578 => (x"ee",x"c0",x"49",x"70"),
  1579 => (x"da",x"c3",x"87",x"d5"),
  1580 => (x"26",x"8e",x"f8",x"87"),
  1581 => (x"20",x"44",x"53",x"4f"),
  1582 => (x"6c",x"69",x"61",x"66"),
  1583 => (x"00",x"2e",x"64",x"65"),
  1584 => (x"74",x"6f",x"6f",x"42"),
  1585 => (x"2e",x"67",x"6e",x"69"),
  1586 => (x"1e",x"00",x"2e",x"2e"),
  1587 => (x"87",x"fa",x"e5",x"c0"),
  1588 => (x"87",x"e9",x"f1",x"c0"),
  1589 => (x"4f",x"26",x"87",x"f6"),
  1590 => (x"c8",x"e8",x"c2",x"1e"),
  1591 => (x"c2",x"78",x"c0",x"48"),
  1592 => (x"c0",x"48",x"f0",x"e7"),
  1593 => (x"87",x"fd",x"fd",x"78"),
  1594 => (x"48",x"c0",x"87",x"e1"),
  1595 => (x"00",x"00",x"4f",x"26"),
  1596 => (x"00",x"00",x"00",x"01"),
  1597 => (x"78",x"45",x"20",x"80"),
  1598 => (x"80",x"00",x"74",x"69"),
  1599 => (x"63",x"61",x"42",x"20"),
  1600 => (x"10",x"25",x"00",x"6b"),
  1601 => (x"2a",x"1c",x"00",x"00"),
  1602 => (x"00",x"00",x"00",x"00"),
  1603 => (x"00",x"10",x"25",x"00"),
  1604 => (x"00",x"2a",x"3a",x"00"),
  1605 => (x"00",x"00",x"00",x"00"),
  1606 => (x"00",x"00",x"10",x"25"),
  1607 => (x"00",x"00",x"2a",x"58"),
  1608 => (x"25",x"00",x"00",x"00"),
  1609 => (x"76",x"00",x"00",x"10"),
  1610 => (x"00",x"00",x"00",x"2a"),
  1611 => (x"10",x"25",x"00",x"00"),
  1612 => (x"2a",x"94",x"00",x"00"),
  1613 => (x"00",x"00",x"00",x"00"),
  1614 => (x"00",x"10",x"25",x"00"),
  1615 => (x"00",x"2a",x"b2",x"00"),
  1616 => (x"00",x"00",x"00",x"00"),
  1617 => (x"00",x"00",x"10",x"25"),
  1618 => (x"00",x"00",x"2a",x"d0"),
  1619 => (x"d8",x"00",x"00",x"00"),
  1620 => (x"00",x"00",x"00",x"10"),
  1621 => (x"00",x"00",x"00",x"00"),
  1622 => (x"13",x"26",x"00",x"00"),
  1623 => (x"00",x"00",x"00",x"00"),
  1624 => (x"00",x"00",x"00",x"00"),
  1625 => (x"00",x"19",x"69",x"00"),
  1626 => (x"4f",x"4f",x"42",x"00"),
  1627 => (x"20",x"20",x"20",x"54"),
  1628 => (x"4d",x"4f",x"52",x"20"),
  1629 => (x"f0",x"fe",x"1e",x"00"),
  1630 => (x"cd",x"78",x"c0",x"48"),
  1631 => (x"26",x"09",x"79",x"09"),
  1632 => (x"fe",x"1e",x"1e",x"4f"),
  1633 => (x"48",x"7e",x"bf",x"f0"),
  1634 => (x"1e",x"4f",x"26",x"26"),
  1635 => (x"c1",x"48",x"f0",x"fe"),
  1636 => (x"1e",x"4f",x"26",x"78"),
  1637 => (x"c0",x"48",x"f0",x"fe"),
  1638 => (x"1e",x"4f",x"26",x"78"),
  1639 => (x"52",x"c0",x"4a",x"71"),
  1640 => (x"0e",x"4f",x"26",x"52"),
  1641 => (x"5d",x"5c",x"5b",x"5e"),
  1642 => (x"71",x"86",x"f4",x"0e"),
  1643 => (x"7e",x"6d",x"97",x"4d"),
  1644 => (x"97",x"4c",x"a5",x"c1"),
  1645 => (x"a6",x"c8",x"48",x"6c"),
  1646 => (x"c4",x"48",x"6e",x"58"),
  1647 => (x"c5",x"05",x"a8",x"66"),
  1648 => (x"c0",x"48",x"ff",x"87"),
  1649 => (x"ca",x"ff",x"87",x"e6"),
  1650 => (x"49",x"a5",x"c2",x"87"),
  1651 => (x"71",x"4b",x"6c",x"97"),
  1652 => (x"6b",x"97",x"4b",x"a3"),
  1653 => (x"7e",x"6c",x"97",x"4b"),
  1654 => (x"80",x"c1",x"48",x"6e"),
  1655 => (x"c7",x"58",x"a6",x"c8"),
  1656 => (x"58",x"a6",x"cc",x"98"),
  1657 => (x"fe",x"7c",x"97",x"70"),
  1658 => (x"48",x"73",x"87",x"e1"),
  1659 => (x"4d",x"26",x"8e",x"f4"),
  1660 => (x"4b",x"26",x"4c",x"26"),
  1661 => (x"5e",x"0e",x"4f",x"26"),
  1662 => (x"f4",x"0e",x"5c",x"5b"),
  1663 => (x"d8",x"4c",x"71",x"86"),
  1664 => (x"ff",x"c3",x"4a",x"66"),
  1665 => (x"4b",x"a4",x"c2",x"9a"),
  1666 => (x"73",x"49",x"6c",x"97"),
  1667 => (x"51",x"72",x"49",x"a1"),
  1668 => (x"6e",x"7e",x"6c",x"97"),
  1669 => (x"c8",x"80",x"c1",x"48"),
  1670 => (x"98",x"c7",x"58",x"a6"),
  1671 => (x"70",x"58",x"a6",x"cc"),
  1672 => (x"ff",x"8e",x"f4",x"54"),
  1673 => (x"1e",x"1e",x"87",x"ca"),
  1674 => (x"e0",x"87",x"e8",x"fd"),
  1675 => (x"c0",x"49",x"4a",x"bf"),
  1676 => (x"02",x"99",x"c0",x"e0"),
  1677 => (x"1e",x"72",x"87",x"cb"),
  1678 => (x"49",x"ee",x"eb",x"c2"),
  1679 => (x"c4",x"87",x"f7",x"fe"),
  1680 => (x"87",x"fd",x"fc",x"86"),
  1681 => (x"c2",x"fd",x"7e",x"70"),
  1682 => (x"4f",x"26",x"26",x"87"),
  1683 => (x"ee",x"eb",x"c2",x"1e"),
  1684 => (x"87",x"c7",x"fd",x"49"),
  1685 => (x"49",x"e6",x"e8",x"c1"),
  1686 => (x"c3",x"87",x"da",x"fc"),
  1687 => (x"4f",x"26",x"87",x"f7"),
  1688 => (x"5c",x"5b",x"5e",x"0e"),
  1689 => (x"4d",x"71",x"0e",x"5d"),
  1690 => (x"49",x"ee",x"eb",x"c2"),
  1691 => (x"70",x"87",x"f4",x"fc"),
  1692 => (x"ab",x"b7",x"c0",x"4b"),
  1693 => (x"87",x"c2",x"c3",x"04"),
  1694 => (x"05",x"ab",x"f0",x"c3"),
  1695 => (x"ed",x"c1",x"87",x"c9"),
  1696 => (x"78",x"c1",x"48",x"c4"),
  1697 => (x"c3",x"87",x"e3",x"c2"),
  1698 => (x"c9",x"05",x"ab",x"e0"),
  1699 => (x"c8",x"ed",x"c1",x"87"),
  1700 => (x"c2",x"78",x"c1",x"48"),
  1701 => (x"ed",x"c1",x"87",x"d4"),
  1702 => (x"c6",x"02",x"bf",x"c8"),
  1703 => (x"a3",x"c0",x"c2",x"87"),
  1704 => (x"73",x"87",x"c2",x"4c"),
  1705 => (x"c4",x"ed",x"c1",x"4c"),
  1706 => (x"e0",x"c0",x"02",x"bf"),
  1707 => (x"c4",x"49",x"74",x"87"),
  1708 => (x"c1",x"91",x"29",x"b7"),
  1709 => (x"74",x"81",x"e4",x"ee"),
  1710 => (x"c2",x"9a",x"cf",x"4a"),
  1711 => (x"72",x"48",x"c1",x"92"),
  1712 => (x"ff",x"4a",x"70",x"30"),
  1713 => (x"69",x"48",x"72",x"ba"),
  1714 => (x"db",x"79",x"70",x"98"),
  1715 => (x"c4",x"49",x"74",x"87"),
  1716 => (x"c1",x"91",x"29",x"b7"),
  1717 => (x"74",x"81",x"e4",x"ee"),
  1718 => (x"c2",x"9a",x"cf",x"4a"),
  1719 => (x"72",x"48",x"c3",x"92"),
  1720 => (x"48",x"4a",x"70",x"30"),
  1721 => (x"79",x"70",x"b0",x"69"),
  1722 => (x"c0",x"05",x"9d",x"75"),
  1723 => (x"d0",x"ff",x"87",x"f0"),
  1724 => (x"78",x"e1",x"c8",x"48"),
  1725 => (x"c5",x"48",x"d4",x"ff"),
  1726 => (x"c8",x"ed",x"c1",x"78"),
  1727 => (x"87",x"c3",x"02",x"bf"),
  1728 => (x"c1",x"78",x"e0",x"c3"),
  1729 => (x"02",x"bf",x"c4",x"ed"),
  1730 => (x"d4",x"ff",x"87",x"c6"),
  1731 => (x"78",x"f0",x"c3",x"48"),
  1732 => (x"7b",x"0b",x"d4",x"ff"),
  1733 => (x"48",x"d0",x"ff",x"0b"),
  1734 => (x"c0",x"78",x"e1",x"c8"),
  1735 => (x"ed",x"c1",x"78",x"e0"),
  1736 => (x"78",x"c0",x"48",x"c8"),
  1737 => (x"48",x"c4",x"ed",x"c1"),
  1738 => (x"eb",x"c2",x"78",x"c0"),
  1739 => (x"f2",x"f9",x"49",x"ee"),
  1740 => (x"c0",x"4b",x"70",x"87"),
  1741 => (x"fc",x"03",x"ab",x"b7"),
  1742 => (x"48",x"c0",x"87",x"fe"),
  1743 => (x"4c",x"26",x"4d",x"26"),
  1744 => (x"4f",x"26",x"4b",x"26"),
  1745 => (x"00",x"00",x"00",x"00"),
  1746 => (x"00",x"00",x"00",x"00"),
  1747 => (x"49",x"4a",x"71",x"1e"),
  1748 => (x"26",x"87",x"cd",x"fc"),
  1749 => (x"4a",x"c0",x"1e",x"4f"),
  1750 => (x"91",x"c4",x"49",x"72"),
  1751 => (x"81",x"e4",x"ee",x"c1"),
  1752 => (x"82",x"c1",x"79",x"c0"),
  1753 => (x"04",x"aa",x"b7",x"d0"),
  1754 => (x"4f",x"26",x"87",x"ee"),
  1755 => (x"5c",x"5b",x"5e",x"0e"),
  1756 => (x"4d",x"71",x"0e",x"5d"),
  1757 => (x"75",x"87",x"dc",x"f8"),
  1758 => (x"2a",x"b7",x"c4",x"4a"),
  1759 => (x"e4",x"ee",x"c1",x"92"),
  1760 => (x"cf",x"4c",x"75",x"82"),
  1761 => (x"6a",x"94",x"c2",x"9c"),
  1762 => (x"2b",x"74",x"4b",x"49"),
  1763 => (x"48",x"c2",x"9b",x"c3"),
  1764 => (x"4c",x"70",x"30",x"74"),
  1765 => (x"48",x"74",x"bc",x"ff"),
  1766 => (x"7a",x"70",x"98",x"71"),
  1767 => (x"73",x"87",x"ec",x"f7"),
  1768 => (x"87",x"d8",x"fe",x"48"),
  1769 => (x"00",x"00",x"00",x"00"),
  1770 => (x"00",x"00",x"00",x"00"),
  1771 => (x"00",x"00",x"00",x"00"),
  1772 => (x"00",x"00",x"00",x"00"),
  1773 => (x"00",x"00",x"00",x"00"),
  1774 => (x"00",x"00",x"00",x"00"),
  1775 => (x"00",x"00",x"00",x"00"),
  1776 => (x"00",x"00",x"00",x"00"),
  1777 => (x"00",x"00",x"00",x"00"),
  1778 => (x"00",x"00",x"00",x"00"),
  1779 => (x"00",x"00",x"00",x"00"),
  1780 => (x"00",x"00",x"00",x"00"),
  1781 => (x"00",x"00",x"00",x"00"),
  1782 => (x"00",x"00",x"00",x"00"),
  1783 => (x"00",x"00",x"00",x"00"),
  1784 => (x"00",x"00",x"00",x"00"),
  1785 => (x"48",x"d0",x"ff",x"1e"),
  1786 => (x"71",x"78",x"e1",x"c8"),
  1787 => (x"08",x"d4",x"ff",x"48"),
  1788 => (x"1e",x"4f",x"26",x"78"),
  1789 => (x"c8",x"48",x"d0",x"ff"),
  1790 => (x"48",x"71",x"78",x"e1"),
  1791 => (x"78",x"08",x"d4",x"ff"),
  1792 => (x"ff",x"48",x"66",x"c4"),
  1793 => (x"26",x"78",x"08",x"d4"),
  1794 => (x"4a",x"71",x"1e",x"4f"),
  1795 => (x"1e",x"49",x"66",x"c4"),
  1796 => (x"de",x"ff",x"49",x"72"),
  1797 => (x"48",x"d0",x"ff",x"87"),
  1798 => (x"26",x"78",x"e0",x"c0"),
  1799 => (x"73",x"1e",x"4f",x"26"),
  1800 => (x"c8",x"4b",x"71",x"1e"),
  1801 => (x"73",x"1e",x"49",x"66"),
  1802 => (x"a2",x"e0",x"c1",x"4a"),
  1803 => (x"87",x"d9",x"ff",x"49"),
  1804 => (x"26",x"87",x"c4",x"26"),
  1805 => (x"26",x"4c",x"26",x"4d"),
  1806 => (x"1e",x"4f",x"26",x"4b"),
  1807 => (x"c3",x"4a",x"d4",x"ff"),
  1808 => (x"d0",x"ff",x"7a",x"ff"),
  1809 => (x"78",x"e1",x"c0",x"48"),
  1810 => (x"eb",x"c2",x"7a",x"de"),
  1811 => (x"49",x"7a",x"bf",x"f8"),
  1812 => (x"70",x"28",x"c8",x"48"),
  1813 => (x"d0",x"48",x"71",x"7a"),
  1814 => (x"71",x"7a",x"70",x"28"),
  1815 => (x"70",x"28",x"d8",x"48"),
  1816 => (x"48",x"d0",x"ff",x"7a"),
  1817 => (x"26",x"78",x"e0",x"c0"),
  1818 => (x"d0",x"ff",x"1e",x"4f"),
  1819 => (x"78",x"c9",x"c8",x"48"),
  1820 => (x"d4",x"ff",x"48",x"71"),
  1821 => (x"4f",x"26",x"78",x"08"),
  1822 => (x"49",x"4a",x"71",x"1e"),
  1823 => (x"d0",x"ff",x"87",x"eb"),
  1824 => (x"26",x"78",x"c8",x"48"),
  1825 => (x"1e",x"73",x"1e",x"4f"),
  1826 => (x"ec",x"c2",x"4b",x"71"),
  1827 => (x"c3",x"02",x"bf",x"c8"),
  1828 => (x"87",x"eb",x"c2",x"87"),
  1829 => (x"c8",x"48",x"d0",x"ff"),
  1830 => (x"48",x"73",x"78",x"c9"),
  1831 => (x"ff",x"b0",x"e0",x"c0"),
  1832 => (x"c2",x"78",x"08",x"d4"),
  1833 => (x"c0",x"48",x"fc",x"eb"),
  1834 => (x"02",x"66",x"c8",x"78"),
  1835 => (x"ff",x"c3",x"87",x"c5"),
  1836 => (x"c0",x"87",x"c2",x"49"),
  1837 => (x"c4",x"ec",x"c2",x"49"),
  1838 => (x"02",x"66",x"cc",x"59"),
  1839 => (x"d5",x"c5",x"87",x"c6"),
  1840 => (x"87",x"c4",x"4a",x"d5"),
  1841 => (x"4a",x"ff",x"ff",x"cf"),
  1842 => (x"5a",x"c8",x"ec",x"c2"),
  1843 => (x"48",x"c8",x"ec",x"c2"),
  1844 => (x"87",x"c4",x"78",x"c1"),
  1845 => (x"4c",x"26",x"4d",x"26"),
  1846 => (x"4f",x"26",x"4b",x"26"),
  1847 => (x"5c",x"5b",x"5e",x"0e"),
  1848 => (x"4a",x"71",x"0e",x"5d"),
  1849 => (x"bf",x"c4",x"ec",x"c2"),
  1850 => (x"02",x"9a",x"72",x"4c"),
  1851 => (x"c8",x"49",x"87",x"cb"),
  1852 => (x"fb",x"f1",x"c1",x"91"),
  1853 => (x"c4",x"83",x"71",x"4b"),
  1854 => (x"fb",x"f5",x"c1",x"87"),
  1855 => (x"13",x"4d",x"c0",x"4b"),
  1856 => (x"c2",x"99",x"74",x"49"),
  1857 => (x"48",x"bf",x"c0",x"ec"),
  1858 => (x"d4",x"ff",x"b8",x"71"),
  1859 => (x"b7",x"c1",x"78",x"08"),
  1860 => (x"b7",x"c8",x"85",x"2c"),
  1861 => (x"87",x"e7",x"04",x"ad"),
  1862 => (x"bf",x"fc",x"eb",x"c2"),
  1863 => (x"c2",x"80",x"c8",x"48"),
  1864 => (x"fe",x"58",x"c0",x"ec"),
  1865 => (x"73",x"1e",x"87",x"ee"),
  1866 => (x"13",x"4b",x"71",x"1e"),
  1867 => (x"cb",x"02",x"9a",x"4a"),
  1868 => (x"fe",x"49",x"72",x"87"),
  1869 => (x"4a",x"13",x"87",x"e6"),
  1870 => (x"87",x"f5",x"05",x"9a"),
  1871 => (x"1e",x"87",x"d9",x"fe"),
  1872 => (x"bf",x"fc",x"eb",x"c2"),
  1873 => (x"fc",x"eb",x"c2",x"49"),
  1874 => (x"78",x"a1",x"c1",x"48"),
  1875 => (x"a9",x"b7",x"c0",x"c4"),
  1876 => (x"ff",x"87",x"db",x"03"),
  1877 => (x"ec",x"c2",x"48",x"d4"),
  1878 => (x"c2",x"78",x"bf",x"c0"),
  1879 => (x"49",x"bf",x"fc",x"eb"),
  1880 => (x"48",x"fc",x"eb",x"c2"),
  1881 => (x"c4",x"78",x"a1",x"c1"),
  1882 => (x"04",x"a9",x"b7",x"c0"),
  1883 => (x"d0",x"ff",x"87",x"e5"),
  1884 => (x"c2",x"78",x"c8",x"48"),
  1885 => (x"c0",x"48",x"c8",x"ec"),
  1886 => (x"00",x"4f",x"26",x"78"),
  1887 => (x"00",x"00",x"00",x"00"),
  1888 => (x"00",x"00",x"00",x"00"),
  1889 => (x"5f",x"5f",x"00",x"00"),
  1890 => (x"00",x"00",x"00",x"00"),
  1891 => (x"03",x"00",x"03",x"03"),
  1892 => (x"14",x"00",x"00",x"03"),
  1893 => (x"7f",x"14",x"7f",x"7f"),
  1894 => (x"00",x"00",x"14",x"7f"),
  1895 => (x"6b",x"6b",x"2e",x"24"),
  1896 => (x"4c",x"00",x"12",x"3a"),
  1897 => (x"6c",x"18",x"36",x"6a"),
  1898 => (x"30",x"00",x"32",x"56"),
  1899 => (x"77",x"59",x"4f",x"7e"),
  1900 => (x"00",x"40",x"68",x"3a"),
  1901 => (x"03",x"07",x"04",x"00"),
  1902 => (x"00",x"00",x"00",x"00"),
  1903 => (x"63",x"3e",x"1c",x"00"),
  1904 => (x"00",x"00",x"00",x"41"),
  1905 => (x"3e",x"63",x"41",x"00"),
  1906 => (x"08",x"00",x"00",x"1c"),
  1907 => (x"1c",x"1c",x"3e",x"2a"),
  1908 => (x"00",x"08",x"2a",x"3e"),
  1909 => (x"3e",x"3e",x"08",x"08"),
  1910 => (x"00",x"00",x"08",x"08"),
  1911 => (x"60",x"e0",x"80",x"00"),
  1912 => (x"00",x"00",x"00",x"00"),
  1913 => (x"08",x"08",x"08",x"08"),
  1914 => (x"00",x"00",x"08",x"08"),
  1915 => (x"60",x"60",x"00",x"00"),
  1916 => (x"40",x"00",x"00",x"00"),
  1917 => (x"0c",x"18",x"30",x"60"),
  1918 => (x"00",x"01",x"03",x"06"),
  1919 => (x"4d",x"59",x"7f",x"3e"),
  1920 => (x"00",x"00",x"3e",x"7f"),
  1921 => (x"7f",x"7f",x"06",x"04"),
  1922 => (x"00",x"00",x"00",x"00"),
  1923 => (x"59",x"71",x"63",x"42"),
  1924 => (x"00",x"00",x"46",x"4f"),
  1925 => (x"49",x"49",x"63",x"22"),
  1926 => (x"18",x"00",x"36",x"7f"),
  1927 => (x"7f",x"13",x"16",x"1c"),
  1928 => (x"00",x"00",x"10",x"7f"),
  1929 => (x"45",x"45",x"67",x"27"),
  1930 => (x"00",x"00",x"39",x"7d"),
  1931 => (x"49",x"4b",x"7e",x"3c"),
  1932 => (x"00",x"00",x"30",x"79"),
  1933 => (x"79",x"71",x"01",x"01"),
  1934 => (x"00",x"00",x"07",x"0f"),
  1935 => (x"49",x"49",x"7f",x"36"),
  1936 => (x"00",x"00",x"36",x"7f"),
  1937 => (x"69",x"49",x"4f",x"06"),
  1938 => (x"00",x"00",x"1e",x"3f"),
  1939 => (x"66",x"66",x"00",x"00"),
  1940 => (x"00",x"00",x"00",x"00"),
  1941 => (x"66",x"e6",x"80",x"00"),
  1942 => (x"00",x"00",x"00",x"00"),
  1943 => (x"14",x"14",x"08",x"08"),
  1944 => (x"00",x"00",x"22",x"22"),
  1945 => (x"14",x"14",x"14",x"14"),
  1946 => (x"00",x"00",x"14",x"14"),
  1947 => (x"14",x"14",x"22",x"22"),
  1948 => (x"00",x"00",x"08",x"08"),
  1949 => (x"59",x"51",x"03",x"02"),
  1950 => (x"3e",x"00",x"06",x"0f"),
  1951 => (x"55",x"5d",x"41",x"7f"),
  1952 => (x"00",x"00",x"1e",x"1f"),
  1953 => (x"09",x"09",x"7f",x"7e"),
  1954 => (x"00",x"00",x"7e",x"7f"),
  1955 => (x"49",x"49",x"7f",x"7f"),
  1956 => (x"00",x"00",x"36",x"7f"),
  1957 => (x"41",x"63",x"3e",x"1c"),
  1958 => (x"00",x"00",x"41",x"41"),
  1959 => (x"63",x"41",x"7f",x"7f"),
  1960 => (x"00",x"00",x"1c",x"3e"),
  1961 => (x"49",x"49",x"7f",x"7f"),
  1962 => (x"00",x"00",x"41",x"41"),
  1963 => (x"09",x"09",x"7f",x"7f"),
  1964 => (x"00",x"00",x"01",x"01"),
  1965 => (x"49",x"41",x"7f",x"3e"),
  1966 => (x"00",x"00",x"7a",x"7b"),
  1967 => (x"08",x"08",x"7f",x"7f"),
  1968 => (x"00",x"00",x"7f",x"7f"),
  1969 => (x"7f",x"7f",x"41",x"00"),
  1970 => (x"00",x"00",x"00",x"41"),
  1971 => (x"40",x"40",x"60",x"20"),
  1972 => (x"7f",x"00",x"3f",x"7f"),
  1973 => (x"36",x"1c",x"08",x"7f"),
  1974 => (x"00",x"00",x"41",x"63"),
  1975 => (x"40",x"40",x"7f",x"7f"),
  1976 => (x"7f",x"00",x"40",x"40"),
  1977 => (x"06",x"0c",x"06",x"7f"),
  1978 => (x"7f",x"00",x"7f",x"7f"),
  1979 => (x"18",x"0c",x"06",x"7f"),
  1980 => (x"00",x"00",x"7f",x"7f"),
  1981 => (x"41",x"41",x"7f",x"3e"),
  1982 => (x"00",x"00",x"3e",x"7f"),
  1983 => (x"09",x"09",x"7f",x"7f"),
  1984 => (x"3e",x"00",x"06",x"0f"),
  1985 => (x"7f",x"61",x"41",x"7f"),
  1986 => (x"00",x"00",x"40",x"7e"),
  1987 => (x"19",x"09",x"7f",x"7f"),
  1988 => (x"00",x"00",x"66",x"7f"),
  1989 => (x"59",x"4d",x"6f",x"26"),
  1990 => (x"00",x"00",x"32",x"7b"),
  1991 => (x"7f",x"7f",x"01",x"01"),
  1992 => (x"00",x"00",x"01",x"01"),
  1993 => (x"40",x"40",x"7f",x"3f"),
  1994 => (x"00",x"00",x"3f",x"7f"),
  1995 => (x"70",x"70",x"3f",x"0f"),
  1996 => (x"7f",x"00",x"0f",x"3f"),
  1997 => (x"30",x"18",x"30",x"7f"),
  1998 => (x"41",x"00",x"7f",x"7f"),
  1999 => (x"1c",x"1c",x"36",x"63"),
  2000 => (x"01",x"41",x"63",x"36"),
  2001 => (x"7c",x"7c",x"06",x"03"),
  2002 => (x"61",x"01",x"03",x"06"),
  2003 => (x"47",x"4d",x"59",x"71"),
  2004 => (x"00",x"00",x"41",x"43"),
  2005 => (x"41",x"7f",x"7f",x"00"),
  2006 => (x"01",x"00",x"00",x"41"),
  2007 => (x"18",x"0c",x"06",x"03"),
  2008 => (x"00",x"40",x"60",x"30"),
  2009 => (x"7f",x"41",x"41",x"00"),
  2010 => (x"08",x"00",x"00",x"7f"),
  2011 => (x"06",x"03",x"06",x"0c"),
  2012 => (x"80",x"00",x"08",x"0c"),
  2013 => (x"80",x"80",x"80",x"80"),
  2014 => (x"00",x"00",x"80",x"80"),
  2015 => (x"07",x"03",x"00",x"00"),
  2016 => (x"00",x"00",x"00",x"04"),
  2017 => (x"54",x"54",x"74",x"20"),
  2018 => (x"00",x"00",x"78",x"7c"),
  2019 => (x"44",x"44",x"7f",x"7f"),
  2020 => (x"00",x"00",x"38",x"7c"),
  2021 => (x"44",x"44",x"7c",x"38"),
  2022 => (x"00",x"00",x"00",x"44"),
  2023 => (x"44",x"44",x"7c",x"38"),
  2024 => (x"00",x"00",x"7f",x"7f"),
  2025 => (x"54",x"54",x"7c",x"38"),
  2026 => (x"00",x"00",x"18",x"5c"),
  2027 => (x"05",x"7f",x"7e",x"04"),
  2028 => (x"00",x"00",x"00",x"05"),
  2029 => (x"a4",x"a4",x"bc",x"18"),
  2030 => (x"00",x"00",x"7c",x"fc"),
  2031 => (x"04",x"04",x"7f",x"7f"),
  2032 => (x"00",x"00",x"78",x"7c"),
  2033 => (x"7d",x"3d",x"00",x"00"),
  2034 => (x"00",x"00",x"00",x"40"),
  2035 => (x"fd",x"80",x"80",x"80"),
  2036 => (x"00",x"00",x"00",x"7d"),
  2037 => (x"38",x"10",x"7f",x"7f"),
  2038 => (x"00",x"00",x"44",x"6c"),
  2039 => (x"7f",x"3f",x"00",x"00"),
  2040 => (x"7c",x"00",x"00",x"40"),
  2041 => (x"0c",x"18",x"0c",x"7c"),
  2042 => (x"00",x"00",x"78",x"7c"),
  2043 => (x"04",x"04",x"7c",x"7c"),
  2044 => (x"00",x"00",x"78",x"7c"),
  2045 => (x"44",x"44",x"7c",x"38"),
  2046 => (x"00",x"00",x"38",x"7c"),
  2047 => (x"24",x"24",x"fc",x"fc"),
  2048 => (x"00",x"00",x"18",x"3c"),
  2049 => (x"24",x"24",x"3c",x"18"),
  2050 => (x"00",x"00",x"fc",x"fc"),
  2051 => (x"04",x"04",x"7c",x"7c"),
  2052 => (x"00",x"00",x"08",x"0c"),
  2053 => (x"54",x"54",x"5c",x"48"),
  2054 => (x"00",x"00",x"20",x"74"),
  2055 => (x"44",x"7f",x"3f",x"04"),
  2056 => (x"00",x"00",x"00",x"44"),
  2057 => (x"40",x"40",x"7c",x"3c"),
  2058 => (x"00",x"00",x"7c",x"7c"),
  2059 => (x"60",x"60",x"3c",x"1c"),
  2060 => (x"3c",x"00",x"1c",x"3c"),
  2061 => (x"60",x"30",x"60",x"7c"),
  2062 => (x"44",x"00",x"3c",x"7c"),
  2063 => (x"38",x"10",x"38",x"6c"),
  2064 => (x"00",x"00",x"44",x"6c"),
  2065 => (x"60",x"e0",x"bc",x"1c"),
  2066 => (x"00",x"00",x"1c",x"3c"),
  2067 => (x"5c",x"74",x"64",x"44"),
  2068 => (x"00",x"00",x"44",x"4c"),
  2069 => (x"77",x"3e",x"08",x"08"),
  2070 => (x"00",x"00",x"41",x"41"),
  2071 => (x"7f",x"7f",x"00",x"00"),
  2072 => (x"00",x"00",x"00",x"00"),
  2073 => (x"3e",x"77",x"41",x"41"),
  2074 => (x"02",x"00",x"08",x"08"),
  2075 => (x"02",x"03",x"01",x"01"),
  2076 => (x"7f",x"00",x"01",x"02"),
  2077 => (x"7f",x"7f",x"7f",x"7f"),
  2078 => (x"08",x"00",x"7f",x"7f"),
  2079 => (x"3e",x"1c",x"1c",x"08"),
  2080 => (x"7f",x"7f",x"7f",x"3e"),
  2081 => (x"1c",x"3e",x"3e",x"7f"),
  2082 => (x"00",x"08",x"08",x"1c"),
  2083 => (x"7c",x"7c",x"18",x"10"),
  2084 => (x"00",x"00",x"10",x"18"),
  2085 => (x"7c",x"7c",x"30",x"10"),
  2086 => (x"10",x"00",x"10",x"30"),
  2087 => (x"78",x"60",x"60",x"30"),
  2088 => (x"42",x"00",x"06",x"1e"),
  2089 => (x"3c",x"18",x"3c",x"66"),
  2090 => (x"78",x"00",x"42",x"66"),
  2091 => (x"c6",x"c2",x"6a",x"38"),
  2092 => (x"60",x"00",x"38",x"6c"),
  2093 => (x"00",x"60",x"00",x"00"),
  2094 => (x"0e",x"00",x"60",x"00"),
  2095 => (x"5d",x"5c",x"5b",x"5e"),
  2096 => (x"4c",x"71",x"1e",x"0e"),
  2097 => (x"bf",x"d9",x"ec",x"c2"),
  2098 => (x"c0",x"4b",x"c0",x"4d"),
  2099 => (x"02",x"ab",x"74",x"1e"),
  2100 => (x"a6",x"c4",x"87",x"c7"),
  2101 => (x"c5",x"78",x"c0",x"48"),
  2102 => (x"48",x"a6",x"c4",x"87"),
  2103 => (x"66",x"c4",x"78",x"c1"),
  2104 => (x"ee",x"49",x"73",x"1e"),
  2105 => (x"86",x"c8",x"87",x"df"),
  2106 => (x"ef",x"49",x"e0",x"c0"),
  2107 => (x"a5",x"c4",x"87",x"ee"),
  2108 => (x"f0",x"49",x"6a",x"4a"),
  2109 => (x"c6",x"f1",x"87",x"f0"),
  2110 => (x"c1",x"85",x"cb",x"87"),
  2111 => (x"ab",x"b7",x"c8",x"83"),
  2112 => (x"87",x"c7",x"ff",x"04"),
  2113 => (x"26",x"4d",x"26",x"26"),
  2114 => (x"26",x"4b",x"26",x"4c"),
  2115 => (x"4a",x"71",x"1e",x"4f"),
  2116 => (x"5a",x"dd",x"ec",x"c2"),
  2117 => (x"48",x"dd",x"ec",x"c2"),
  2118 => (x"fe",x"49",x"78",x"c7"),
  2119 => (x"4f",x"26",x"87",x"dd"),
  2120 => (x"71",x"1e",x"73",x"1e"),
  2121 => (x"aa",x"b7",x"c0",x"4a"),
  2122 => (x"c2",x"87",x"d3",x"03"),
  2123 => (x"05",x"bf",x"dc",x"d2"),
  2124 => (x"4b",x"c1",x"87",x"c4"),
  2125 => (x"4b",x"c0",x"87",x"c2"),
  2126 => (x"5b",x"e0",x"d2",x"c2"),
  2127 => (x"d2",x"c2",x"87",x"c4"),
  2128 => (x"d2",x"c2",x"5a",x"e0"),
  2129 => (x"c1",x"4a",x"bf",x"dc"),
  2130 => (x"a2",x"c0",x"c1",x"9a"),
  2131 => (x"87",x"e8",x"ec",x"49"),
  2132 => (x"d2",x"c2",x"48",x"fc"),
  2133 => (x"fe",x"78",x"bf",x"dc"),
  2134 => (x"71",x"1e",x"87",x"ef"),
  2135 => (x"1e",x"66",x"c4",x"4a"),
  2136 => (x"f9",x"ea",x"49",x"72"),
  2137 => (x"4f",x"26",x"26",x"87"),
  2138 => (x"48",x"d4",x"ff",x"1e"),
  2139 => (x"ff",x"78",x"ff",x"c3"),
  2140 => (x"e1",x"c0",x"48",x"d0"),
  2141 => (x"48",x"d4",x"ff",x"78"),
  2142 => (x"48",x"71",x"78",x"c1"),
  2143 => (x"d4",x"ff",x"30",x"c4"),
  2144 => (x"d0",x"ff",x"78",x"08"),
  2145 => (x"78",x"e0",x"c0",x"48"),
  2146 => (x"c2",x"1e",x"4f",x"26"),
  2147 => (x"49",x"bf",x"dc",x"d2"),
  2148 => (x"c2",x"87",x"f9",x"e6"),
  2149 => (x"e8",x"48",x"d1",x"ec"),
  2150 => (x"ec",x"c2",x"78",x"bf"),
  2151 => (x"bf",x"ec",x"48",x"cd"),
  2152 => (x"d1",x"ec",x"c2",x"78"),
  2153 => (x"c3",x"49",x"4a",x"bf"),
  2154 => (x"b7",x"c8",x"99",x"ff"),
  2155 => (x"71",x"48",x"72",x"2a"),
  2156 => (x"d9",x"ec",x"c2",x"b0"),
  2157 => (x"0e",x"4f",x"26",x"58"),
  2158 => (x"5d",x"5c",x"5b",x"5e"),
  2159 => (x"ff",x"4b",x"71",x"0e"),
  2160 => (x"ec",x"c2",x"87",x"c8"),
  2161 => (x"50",x"c0",x"48",x"cc"),
  2162 => (x"df",x"e6",x"49",x"73"),
  2163 => (x"4c",x"49",x"70",x"87"),
  2164 => (x"ee",x"cb",x"9c",x"c2"),
  2165 => (x"87",x"cc",x"cb",x"49"),
  2166 => (x"ec",x"c2",x"4d",x"70"),
  2167 => (x"05",x"bf",x"97",x"cc"),
  2168 => (x"d0",x"87",x"e2",x"c1"),
  2169 => (x"ec",x"c2",x"49",x"66"),
  2170 => (x"05",x"99",x"bf",x"d5"),
  2171 => (x"66",x"d4",x"87",x"d6"),
  2172 => (x"cd",x"ec",x"c2",x"49"),
  2173 => (x"cb",x"05",x"99",x"bf"),
  2174 => (x"e5",x"49",x"73",x"87"),
  2175 => (x"98",x"70",x"87",x"ee"),
  2176 => (x"87",x"c1",x"c1",x"02"),
  2177 => (x"c1",x"fe",x"4c",x"c1"),
  2178 => (x"ca",x"49",x"75",x"87"),
  2179 => (x"98",x"70",x"87",x"e2"),
  2180 => (x"c2",x"87",x"c6",x"02"),
  2181 => (x"c1",x"48",x"cc",x"ec"),
  2182 => (x"cc",x"ec",x"c2",x"50"),
  2183 => (x"c0",x"05",x"bf",x"97"),
  2184 => (x"ec",x"c2",x"87",x"e3"),
  2185 => (x"d0",x"49",x"bf",x"d5"),
  2186 => (x"ff",x"05",x"99",x"66"),
  2187 => (x"ec",x"c2",x"87",x"d6"),
  2188 => (x"d4",x"49",x"bf",x"cd"),
  2189 => (x"ff",x"05",x"99",x"66"),
  2190 => (x"49",x"73",x"87",x"ca"),
  2191 => (x"70",x"87",x"ed",x"e4"),
  2192 => (x"ff",x"fe",x"05",x"98"),
  2193 => (x"fa",x"48",x"74",x"87"),
  2194 => (x"5e",x"0e",x"87",x"fb"),
  2195 => (x"0e",x"5d",x"5c",x"5b"),
  2196 => (x"4d",x"c0",x"86",x"f8"),
  2197 => (x"7e",x"bf",x"ec",x"4c"),
  2198 => (x"c2",x"48",x"a6",x"c4"),
  2199 => (x"78",x"bf",x"d9",x"ec"),
  2200 => (x"1e",x"c0",x"1e",x"c1"),
  2201 => (x"ce",x"fd",x"49",x"c7"),
  2202 => (x"70",x"86",x"c8",x"87"),
  2203 => (x"87",x"cd",x"02",x"98"),
  2204 => (x"eb",x"fa",x"49",x"ff"),
  2205 => (x"49",x"da",x"c1",x"87"),
  2206 => (x"c1",x"87",x"f1",x"e3"),
  2207 => (x"cc",x"ec",x"c2",x"4d"),
  2208 => (x"cf",x"02",x"bf",x"97"),
  2209 => (x"d4",x"d2",x"c2",x"87"),
  2210 => (x"b9",x"c1",x"49",x"bf"),
  2211 => (x"59",x"d8",x"d2",x"c2"),
  2212 => (x"87",x"d4",x"fb",x"71"),
  2213 => (x"bf",x"d1",x"ec",x"c2"),
  2214 => (x"dc",x"d2",x"c2",x"4b"),
  2215 => (x"e9",x"c0",x"05",x"bf"),
  2216 => (x"49",x"fd",x"c3",x"87"),
  2217 => (x"c3",x"87",x"c5",x"e3"),
  2218 => (x"ff",x"e2",x"49",x"fa"),
  2219 => (x"c3",x"49",x"73",x"87"),
  2220 => (x"1e",x"71",x"99",x"ff"),
  2221 => (x"e1",x"fa",x"49",x"c0"),
  2222 => (x"c8",x"49",x"73",x"87"),
  2223 => (x"1e",x"71",x"29",x"b7"),
  2224 => (x"d5",x"fa",x"49",x"c1"),
  2225 => (x"c5",x"86",x"c8",x"87"),
  2226 => (x"ec",x"c2",x"87",x"f4"),
  2227 => (x"9b",x"4b",x"bf",x"d5"),
  2228 => (x"c2",x"87",x"dd",x"02"),
  2229 => (x"49",x"bf",x"d8",x"d2"),
  2230 => (x"70",x"87",x"d5",x"c7"),
  2231 => (x"87",x"c4",x"05",x"98"),
  2232 => (x"87",x"d2",x"4b",x"c0"),
  2233 => (x"c6",x"49",x"e0",x"c2"),
  2234 => (x"d2",x"c2",x"87",x"fa"),
  2235 => (x"87",x"c6",x"58",x"dc"),
  2236 => (x"48",x"d8",x"d2",x"c2"),
  2237 => (x"49",x"73",x"78",x"c0"),
  2238 => (x"cd",x"05",x"99",x"c2"),
  2239 => (x"49",x"eb",x"c3",x"87"),
  2240 => (x"70",x"87",x"e9",x"e1"),
  2241 => (x"02",x"99",x"c2",x"49"),
  2242 => (x"4c",x"fb",x"87",x"c2"),
  2243 => (x"99",x"c1",x"49",x"73"),
  2244 => (x"c3",x"87",x"cd",x"05"),
  2245 => (x"d3",x"e1",x"49",x"f4"),
  2246 => (x"c2",x"49",x"70",x"87"),
  2247 => (x"87",x"c2",x"02",x"99"),
  2248 => (x"49",x"73",x"4c",x"fa"),
  2249 => (x"cd",x"05",x"99",x"c8"),
  2250 => (x"49",x"f5",x"c3",x"87"),
  2251 => (x"70",x"87",x"fd",x"e0"),
  2252 => (x"02",x"99",x"c2",x"49"),
  2253 => (x"ec",x"c2",x"87",x"d5"),
  2254 => (x"ca",x"02",x"bf",x"dd"),
  2255 => (x"88",x"c1",x"48",x"87"),
  2256 => (x"58",x"e1",x"ec",x"c2"),
  2257 => (x"ff",x"87",x"c2",x"c0"),
  2258 => (x"73",x"4d",x"c1",x"4c"),
  2259 => (x"05",x"99",x"c4",x"49"),
  2260 => (x"f2",x"c3",x"87",x"cd"),
  2261 => (x"87",x"d4",x"e0",x"49"),
  2262 => (x"99",x"c2",x"49",x"70"),
  2263 => (x"c2",x"87",x"dc",x"02"),
  2264 => (x"7e",x"bf",x"dd",x"ec"),
  2265 => (x"a8",x"b7",x"c7",x"48"),
  2266 => (x"87",x"cb",x"c0",x"03"),
  2267 => (x"80",x"c1",x"48",x"6e"),
  2268 => (x"58",x"e1",x"ec",x"c2"),
  2269 => (x"fe",x"87",x"c2",x"c0"),
  2270 => (x"c3",x"4d",x"c1",x"4c"),
  2271 => (x"df",x"ff",x"49",x"fd"),
  2272 => (x"49",x"70",x"87",x"ea"),
  2273 => (x"d5",x"02",x"99",x"c2"),
  2274 => (x"dd",x"ec",x"c2",x"87"),
  2275 => (x"c9",x"c0",x"02",x"bf"),
  2276 => (x"dd",x"ec",x"c2",x"87"),
  2277 => (x"c0",x"78",x"c0",x"48"),
  2278 => (x"4c",x"fd",x"87",x"c2"),
  2279 => (x"fa",x"c3",x"4d",x"c1"),
  2280 => (x"c7",x"df",x"ff",x"49"),
  2281 => (x"c2",x"49",x"70",x"87"),
  2282 => (x"d9",x"c0",x"02",x"99"),
  2283 => (x"dd",x"ec",x"c2",x"87"),
  2284 => (x"b7",x"c7",x"48",x"bf"),
  2285 => (x"c9",x"c0",x"03",x"a8"),
  2286 => (x"dd",x"ec",x"c2",x"87"),
  2287 => (x"c0",x"78",x"c7",x"48"),
  2288 => (x"4c",x"fc",x"87",x"c2"),
  2289 => (x"b7",x"c0",x"4d",x"c1"),
  2290 => (x"d3",x"c0",x"03",x"ac"),
  2291 => (x"48",x"66",x"c4",x"87"),
  2292 => (x"70",x"80",x"d8",x"c1"),
  2293 => (x"02",x"bf",x"6e",x"7e"),
  2294 => (x"4b",x"87",x"c5",x"c0"),
  2295 => (x"0f",x"73",x"49",x"74"),
  2296 => (x"f0",x"c3",x"1e",x"c0"),
  2297 => (x"49",x"da",x"c1",x"1e"),
  2298 => (x"c8",x"87",x"cc",x"f7"),
  2299 => (x"02",x"98",x"70",x"86"),
  2300 => (x"c2",x"87",x"d8",x"c0"),
  2301 => (x"7e",x"bf",x"dd",x"ec"),
  2302 => (x"91",x"cb",x"49",x"6e"),
  2303 => (x"71",x"4a",x"66",x"c4"),
  2304 => (x"c0",x"02",x"6a",x"82"),
  2305 => (x"6e",x"4b",x"87",x"c5"),
  2306 => (x"75",x"0f",x"73",x"49"),
  2307 => (x"c8",x"c0",x"02",x"9d"),
  2308 => (x"dd",x"ec",x"c2",x"87"),
  2309 => (x"e2",x"f2",x"49",x"bf"),
  2310 => (x"e0",x"d2",x"c2",x"87"),
  2311 => (x"dd",x"c0",x"02",x"bf"),
  2312 => (x"cb",x"c2",x"49",x"87"),
  2313 => (x"02",x"98",x"70",x"87"),
  2314 => (x"c2",x"87",x"d3",x"c0"),
  2315 => (x"49",x"bf",x"dd",x"ec"),
  2316 => (x"c0",x"87",x"c8",x"f2"),
  2317 => (x"87",x"e8",x"f3",x"49"),
  2318 => (x"48",x"e0",x"d2",x"c2"),
  2319 => (x"8e",x"f8",x"78",x"c0"),
  2320 => (x"0e",x"87",x"c2",x"f3"),
  2321 => (x"5d",x"5c",x"5b",x"5e"),
  2322 => (x"4c",x"71",x"1e",x"0e"),
  2323 => (x"bf",x"d9",x"ec",x"c2"),
  2324 => (x"a1",x"cd",x"c1",x"49"),
  2325 => (x"81",x"d1",x"c1",x"4d"),
  2326 => (x"9c",x"74",x"7e",x"69"),
  2327 => (x"c4",x"87",x"cf",x"02"),
  2328 => (x"7b",x"74",x"4b",x"a5"),
  2329 => (x"bf",x"d9",x"ec",x"c2"),
  2330 => (x"87",x"e1",x"f2",x"49"),
  2331 => (x"9c",x"74",x"7b",x"6e"),
  2332 => (x"c0",x"87",x"c4",x"05"),
  2333 => (x"c1",x"87",x"c2",x"4b"),
  2334 => (x"f2",x"49",x"73",x"4b"),
  2335 => (x"66",x"d4",x"87",x"e2"),
  2336 => (x"49",x"87",x"c7",x"02"),
  2337 => (x"4a",x"70",x"87",x"de"),
  2338 => (x"4a",x"c0",x"87",x"c2"),
  2339 => (x"5a",x"e4",x"d2",x"c2"),
  2340 => (x"87",x"f1",x"f1",x"26"),
  2341 => (x"00",x"00",x"00",x"00"),
  2342 => (x"00",x"00",x"00",x"00"),
  2343 => (x"00",x"00",x"00",x"00"),
  2344 => (x"00",x"00",x"00",x"00"),
  2345 => (x"ff",x"4a",x"71",x"1e"),
  2346 => (x"72",x"49",x"bf",x"c8"),
  2347 => (x"4f",x"26",x"48",x"a1"),
  2348 => (x"bf",x"c8",x"ff",x"1e"),
  2349 => (x"c0",x"c0",x"fe",x"89"),
  2350 => (x"a9",x"c0",x"c0",x"c0"),
  2351 => (x"c0",x"87",x"c4",x"01"),
  2352 => (x"c1",x"87",x"c2",x"4a"),
  2353 => (x"26",x"48",x"72",x"4a"),
  2354 => (x"5b",x"5e",x"0e",x"4f"),
  2355 => (x"71",x"0e",x"5d",x"5c"),
  2356 => (x"4c",x"d4",x"ff",x"4b"),
  2357 => (x"c0",x"48",x"66",x"d0"),
  2358 => (x"ff",x"49",x"d6",x"78"),
  2359 => (x"c3",x"87",x"c5",x"dc"),
  2360 => (x"49",x"6c",x"7c",x"ff"),
  2361 => (x"71",x"99",x"ff",x"c3"),
  2362 => (x"f0",x"c3",x"49",x"4d"),
  2363 => (x"a9",x"e0",x"c1",x"99"),
  2364 => (x"c3",x"87",x"cb",x"05"),
  2365 => (x"48",x"6c",x"7c",x"ff"),
  2366 => (x"66",x"d0",x"98",x"c3"),
  2367 => (x"ff",x"c3",x"78",x"08"),
  2368 => (x"49",x"4a",x"6c",x"7c"),
  2369 => (x"ff",x"c3",x"31",x"c8"),
  2370 => (x"71",x"4a",x"6c",x"7c"),
  2371 => (x"c8",x"49",x"72",x"b2"),
  2372 => (x"7c",x"ff",x"c3",x"31"),
  2373 => (x"b2",x"71",x"4a",x"6c"),
  2374 => (x"31",x"c8",x"49",x"72"),
  2375 => (x"6c",x"7c",x"ff",x"c3"),
  2376 => (x"ff",x"b2",x"71",x"4a"),
  2377 => (x"e0",x"c0",x"48",x"d0"),
  2378 => (x"02",x"9b",x"73",x"78"),
  2379 => (x"7b",x"72",x"87",x"c2"),
  2380 => (x"4d",x"26",x"48",x"75"),
  2381 => (x"4b",x"26",x"4c",x"26"),
  2382 => (x"26",x"1e",x"4f",x"26"),
  2383 => (x"5b",x"5e",x"0e",x"4f"),
  2384 => (x"86",x"f8",x"0e",x"5c"),
  2385 => (x"a6",x"c8",x"1e",x"76"),
  2386 => (x"87",x"fd",x"fd",x"49"),
  2387 => (x"4b",x"70",x"86",x"c4"),
  2388 => (x"a8",x"c8",x"48",x"6e"),
  2389 => (x"87",x"f0",x"c2",x"03"),
  2390 => (x"f0",x"c3",x"4a",x"73"),
  2391 => (x"aa",x"d0",x"c1",x"9a"),
  2392 => (x"c1",x"87",x"c7",x"02"),
  2393 => (x"c2",x"05",x"aa",x"e0"),
  2394 => (x"49",x"73",x"87",x"de"),
  2395 => (x"c3",x"02",x"99",x"c8"),
  2396 => (x"87",x"c6",x"ff",x"87"),
  2397 => (x"9c",x"c3",x"4c",x"73"),
  2398 => (x"c1",x"05",x"ac",x"c2"),
  2399 => (x"66",x"c4",x"87",x"c2"),
  2400 => (x"71",x"31",x"c9",x"49"),
  2401 => (x"4a",x"66",x"c4",x"1e"),
  2402 => (x"ec",x"c2",x"92",x"d4"),
  2403 => (x"81",x"72",x"49",x"e1"),
  2404 => (x"87",x"f3",x"d0",x"fe"),
  2405 => (x"d9",x"ff",x"49",x"d8"),
  2406 => (x"c0",x"c8",x"87",x"ca"),
  2407 => (x"fe",x"da",x"c2",x"1e"),
  2408 => (x"f9",x"ec",x"fd",x"49"),
  2409 => (x"48",x"d0",x"ff",x"87"),
  2410 => (x"c2",x"78",x"e0",x"c0"),
  2411 => (x"cc",x"1e",x"fe",x"da"),
  2412 => (x"92",x"d4",x"4a",x"66"),
  2413 => (x"49",x"e1",x"ec",x"c2"),
  2414 => (x"ce",x"fe",x"81",x"72"),
  2415 => (x"86",x"cc",x"87",x"fb"),
  2416 => (x"c1",x"05",x"ac",x"c1"),
  2417 => (x"66",x"c4",x"87",x"c2"),
  2418 => (x"71",x"31",x"c9",x"49"),
  2419 => (x"4a",x"66",x"c4",x"1e"),
  2420 => (x"ec",x"c2",x"92",x"d4"),
  2421 => (x"81",x"72",x"49",x"e1"),
  2422 => (x"87",x"eb",x"cf",x"fe"),
  2423 => (x"1e",x"fe",x"da",x"c2"),
  2424 => (x"d4",x"4a",x"66",x"c8"),
  2425 => (x"e1",x"ec",x"c2",x"92"),
  2426 => (x"fe",x"81",x"72",x"49"),
  2427 => (x"d7",x"87",x"fc",x"cc"),
  2428 => (x"ef",x"d7",x"ff",x"49"),
  2429 => (x"1e",x"c0",x"c8",x"87"),
  2430 => (x"49",x"fe",x"da",x"c2"),
  2431 => (x"87",x"f7",x"ea",x"fd"),
  2432 => (x"d0",x"ff",x"86",x"cc"),
  2433 => (x"78",x"e0",x"c0",x"48"),
  2434 => (x"e7",x"fc",x"8e",x"f8"),
  2435 => (x"5b",x"5e",x"0e",x"87"),
  2436 => (x"1e",x"0e",x"5d",x"5c"),
  2437 => (x"d4",x"ff",x"4d",x"71"),
  2438 => (x"7e",x"66",x"d4",x"4c"),
  2439 => (x"a8",x"b7",x"c3",x"48"),
  2440 => (x"c0",x"87",x"c5",x"06"),
  2441 => (x"87",x"e9",x"c1",x"48"),
  2442 => (x"dd",x"fe",x"49",x"75"),
  2443 => (x"1e",x"75",x"87",x"e0"),
  2444 => (x"d4",x"4b",x"66",x"c4"),
  2445 => (x"e1",x"ec",x"c2",x"93"),
  2446 => (x"fe",x"49",x"73",x"83"),
  2447 => (x"c8",x"87",x"fa",x"c6"),
  2448 => (x"ff",x"4b",x"6b",x"83"),
  2449 => (x"e1",x"c8",x"48",x"d0"),
  2450 => (x"73",x"7c",x"dd",x"78"),
  2451 => (x"98",x"ff",x"c3",x"48"),
  2452 => (x"49",x"73",x"7c",x"70"),
  2453 => (x"71",x"29",x"b7",x"c8"),
  2454 => (x"98",x"ff",x"c3",x"48"),
  2455 => (x"49",x"73",x"7c",x"70"),
  2456 => (x"71",x"29",x"b7",x"d0"),
  2457 => (x"98",x"ff",x"c3",x"48"),
  2458 => (x"48",x"73",x"7c",x"70"),
  2459 => (x"70",x"28",x"b7",x"d8"),
  2460 => (x"7c",x"7c",x"c0",x"7c"),
  2461 => (x"7c",x"7c",x"7c",x"7c"),
  2462 => (x"7c",x"7c",x"7c",x"7c"),
  2463 => (x"d0",x"ff",x"7c",x"7c"),
  2464 => (x"78",x"e0",x"c0",x"48"),
  2465 => (x"dc",x"1e",x"66",x"c4"),
  2466 => (x"fc",x"d5",x"ff",x"49"),
  2467 => (x"73",x"86",x"c8",x"87"),
  2468 => (x"dd",x"fa",x"26",x"48"),
  2469 => (x"dd",x"fa",x"26",x"87"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

